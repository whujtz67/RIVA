package vlsu_shuffle_pkg;

  // Input sequential index, output shuffle index
  // Used in Deshuffle Unit to convert sequential index to shuffle index
  function automatic logic [{$clog2(riva_pkg::DLEN*riva_pkg::MaxNrLanes/4)}-1:0] query_shf_idx(input int NrLanes, input int seqNbIdx, input riscv_mv_pkg::vew_e ew);
    // Lookup tables for each lane configuration
    automatic logic [5-1:0] lut_1lane [0:31][0:3] = '{
      '{5'd000, 5'd000, 5'd000, 5'd000}, '{5'd008, 5'd001, 5'd001, 5'd001}, '{5'd016, 5'd008, 5'd002, 5'd002}, '{5'd024, 5'd009, 5'd003, 5'd003},
      '{5'd004, 5'd016, 5'd008, 5'd004}, '{5'd012, 5'd017, 5'd009, 5'd005}, '{5'd020, 5'd024, 5'd010, 5'd006}, '{5'd028, 5'd025, 5'd011, 5'd007},
      '{5'd002, 5'd004, 5'd016, 5'd008}, '{5'd010, 5'd005, 5'd017, 5'd009}, '{5'd018, 5'd012, 5'd018, 5'd010}, '{5'd026, 5'd013, 5'd019, 5'd011},
      '{5'd006, 5'd020, 5'd024, 5'd012}, '{5'd014, 5'd021, 5'd025, 5'd013}, '{5'd022, 5'd028, 5'd026, 5'd014}, '{5'd030, 5'd029, 5'd027, 5'd015},
      '{5'd001, 5'd002, 5'd004, 5'd016}, '{5'd009, 5'd003, 5'd005, 5'd017}, '{5'd017, 5'd010, 5'd006, 5'd018}, '{5'd025, 5'd011, 5'd007, 5'd019},
      '{5'd005, 5'd018, 5'd012, 5'd020}, '{5'd013, 5'd019, 5'd013, 5'd021}, '{5'd021, 5'd026, 5'd014, 5'd022}, '{5'd029, 5'd027, 5'd015, 5'd023},
      '{5'd003, 5'd006, 5'd020, 5'd024}, '{5'd011, 5'd007, 5'd021, 5'd025}, '{5'd019, 5'd014, 5'd022, 5'd026}, '{5'd027, 5'd015, 5'd023, 5'd027},
      '{5'd007, 5'd022, 5'd028, 5'd028}, '{5'd015, 5'd023, 5'd029, 5'd029}, '{5'd023, 5'd030, 5'd030, 5'd030}, '{5'd031, 5'd031, 5'd031, 5'd031}
    };
    automatic logic [6-1:0] lut_2lane [0:63][0:3] = '{
      '{6'd000, 6'd000, 6'd000, 6'd000}, '{6'd032, 6'd001, 6'd001, 6'd001}, '{6'd008, 6'd032, 6'd002, 6'd002}, '{6'd040, 6'd033, 6'd003, 6'd003},
      '{6'd016, 6'd008, 6'd032, 6'd004}, '{6'd048, 6'd009, 6'd033, 6'd005}, '{6'd024, 6'd040, 6'd034, 6'd006}, '{6'd056, 6'd041, 6'd035, 6'd007},
      '{6'd004, 6'd016, 6'd008, 6'd032}, '{6'd036, 6'd017, 6'd009, 6'd033}, '{6'd012, 6'd048, 6'd010, 6'd034}, '{6'd044, 6'd049, 6'd011, 6'd035},
      '{6'd020, 6'd024, 6'd040, 6'd036}, '{6'd052, 6'd025, 6'd041, 6'd037}, '{6'd028, 6'd056, 6'd042, 6'd038}, '{6'd060, 6'd057, 6'd043, 6'd039},
      '{6'd002, 6'd004, 6'd016, 6'd008}, '{6'd034, 6'd005, 6'd017, 6'd009}, '{6'd010, 6'd036, 6'd018, 6'd010}, '{6'd042, 6'd037, 6'd019, 6'd011},
      '{6'd018, 6'd012, 6'd048, 6'd012}, '{6'd050, 6'd013, 6'd049, 6'd013}, '{6'd026, 6'd044, 6'd050, 6'd014}, '{6'd058, 6'd045, 6'd051, 6'd015},
      '{6'd006, 6'd020, 6'd024, 6'd040}, '{6'd038, 6'd021, 6'd025, 6'd041}, '{6'd014, 6'd052, 6'd026, 6'd042}, '{6'd046, 6'd053, 6'd027, 6'd043},
      '{6'd022, 6'd028, 6'd056, 6'd044}, '{6'd054, 6'd029, 6'd057, 6'd045}, '{6'd030, 6'd060, 6'd058, 6'd046}, '{6'd062, 6'd061, 6'd059, 6'd047},
      '{6'd001, 6'd002, 6'd004, 6'd016}, '{6'd033, 6'd003, 6'd005, 6'd017}, '{6'd009, 6'd034, 6'd006, 6'd018}, '{6'd041, 6'd035, 6'd007, 6'd019},
      '{6'd017, 6'd010, 6'd036, 6'd020}, '{6'd049, 6'd011, 6'd037, 6'd021}, '{6'd025, 6'd042, 6'd038, 6'd022}, '{6'd057, 6'd043, 6'd039, 6'd023},
      '{6'd005, 6'd018, 6'd012, 6'd048}, '{6'd037, 6'd019, 6'd013, 6'd049}, '{6'd013, 6'd050, 6'd014, 6'd050}, '{6'd045, 6'd051, 6'd015, 6'd051},
      '{6'd021, 6'd026, 6'd044, 6'd052}, '{6'd053, 6'd027, 6'd045, 6'd053}, '{6'd029, 6'd058, 6'd046, 6'd054}, '{6'd061, 6'd059, 6'd047, 6'd055},
      '{6'd003, 6'd006, 6'd020, 6'd024}, '{6'd035, 6'd007, 6'd021, 6'd025}, '{6'd011, 6'd038, 6'd022, 6'd026}, '{6'd043, 6'd039, 6'd023, 6'd027},
      '{6'd019, 6'd014, 6'd052, 6'd028}, '{6'd051, 6'd015, 6'd053, 6'd029}, '{6'd027, 6'd046, 6'd054, 6'd030}, '{6'd059, 6'd047, 6'd055, 6'd031},
      '{6'd007, 6'd022, 6'd028, 6'd056}, '{6'd039, 6'd023, 6'd029, 6'd057}, '{6'd015, 6'd054, 6'd030, 6'd058}, '{6'd047, 6'd055, 6'd031, 6'd059},
      '{6'd023, 6'd030, 6'd060, 6'd060}, '{6'd055, 6'd031, 6'd061, 6'd061}, '{6'd031, 6'd062, 6'd062, 6'd062}, '{6'd063, 6'd063, 6'd063, 6'd063}
    };
    automatic logic [7-1:0] lut_4lane [0:127][0:3] = '{
      '{7'd000, 7'd000, 7'd000, 7'd000}, '{7'd032, 7'd001, 7'd001, 7'd001}, '{7'd064, 7'd032, 7'd002, 7'd002}, '{7'd096, 7'd033, 7'd003, 7'd003},
      '{7'd016, 7'd008, 7'd032, 7'd004}, '{7'd048, 7'd009, 7'd033, 7'd005}, '{7'd080, 7'd040, 7'd034, 7'd006}, '{7'd112, 7'd041, 7'd035, 7'd007},
      '{7'd004, 7'd016, 7'd008, 7'd032}, '{7'd036, 7'd017, 7'd009, 7'd033}, '{7'd068, 7'd048, 7'd010, 7'd034}, '{7'd100, 7'd049, 7'd011, 7'd035},
      '{7'd020, 7'd024, 7'd040, 7'd036}, '{7'd052, 7'd025, 7'd041, 7'd037}, '{7'd084, 7'd056, 7'd042, 7'd038}, '{7'd116, 7'd057, 7'd043, 7'd039},
      '{7'd002, 7'd004, 7'd016, 7'd008}, '{7'd034, 7'd005, 7'd017, 7'd009}, '{7'd066, 7'd036, 7'd018, 7'd010}, '{7'd098, 7'd037, 7'd019, 7'd011},
      '{7'd018, 7'd012, 7'd048, 7'd012}, '{7'd050, 7'd013, 7'd049, 7'd013}, '{7'd082, 7'd044, 7'd050, 7'd014}, '{7'd114, 7'd045, 7'd051, 7'd015},
      '{7'd006, 7'd020, 7'd024, 7'd040}, '{7'd038, 7'd021, 7'd025, 7'd041}, '{7'd070, 7'd052, 7'd026, 7'd042}, '{7'd102, 7'd053, 7'd027, 7'd043},
      '{7'd022, 7'd028, 7'd056, 7'd044}, '{7'd054, 7'd029, 7'd057, 7'd045}, '{7'd086, 7'd060, 7'd058, 7'd046}, '{7'd118, 7'd061, 7'd059, 7'd047},
      '{7'd001, 7'd002, 7'd004, 7'd016}, '{7'd033, 7'd003, 7'd005, 7'd017}, '{7'd065, 7'd034, 7'd006, 7'd018}, '{7'd097, 7'd035, 7'd007, 7'd019},
      '{7'd017, 7'd010, 7'd036, 7'd020}, '{7'd049, 7'd011, 7'd037, 7'd021}, '{7'd081, 7'd042, 7'd038, 7'd022}, '{7'd113, 7'd043, 7'd039, 7'd023},
      '{7'd005, 7'd018, 7'd012, 7'd048}, '{7'd037, 7'd019, 7'd013, 7'd049}, '{7'd069, 7'd050, 7'd014, 7'd050}, '{7'd101, 7'd051, 7'd015, 7'd051},
      '{7'd021, 7'd026, 7'd044, 7'd052}, '{7'd053, 7'd027, 7'd045, 7'd053}, '{7'd085, 7'd058, 7'd046, 7'd054}, '{7'd117, 7'd059, 7'd047, 7'd055},
      '{7'd003, 7'd006, 7'd020, 7'd024}, '{7'd035, 7'd007, 7'd021, 7'd025}, '{7'd067, 7'd038, 7'd022, 7'd026}, '{7'd099, 7'd039, 7'd023, 7'd027},
      '{7'd019, 7'd014, 7'd052, 7'd028}, '{7'd051, 7'd015, 7'd053, 7'd029}, '{7'd083, 7'd046, 7'd054, 7'd030}, '{7'd115, 7'd047, 7'd055, 7'd031},
      '{7'd007, 7'd022, 7'd028, 7'd056}, '{7'd039, 7'd023, 7'd029, 7'd057}, '{7'd071, 7'd054, 7'd030, 7'd058}, '{7'd103, 7'd055, 7'd031, 7'd059},
      '{7'd023, 7'd030, 7'd060, 7'd060}, '{7'd055, 7'd031, 7'd061, 7'd061}, '{7'd087, 7'd062, 7'd062, 7'd062}, '{7'd119, 7'd063, 7'd063, 7'd063},
      '{7'd008, 7'd064, 7'd096, 7'd064}, '{7'd040, 7'd065, 7'd097, 7'd065}, '{7'd072, 7'd096, 7'd098, 7'd066}, '{7'd104, 7'd097, 7'd099, 7'd067},
      '{7'd024, 7'd072, 7'd100, 7'd068}, '{7'd056, 7'd073, 7'd101, 7'd069}, '{7'd088, 7'd104, 7'd102, 7'd070}, '{7'd120, 7'd105, 7'd103, 7'd071},
      '{7'd012, 7'd080, 7'd104, 7'd072}, '{7'd044, 7'd081, 7'd105, 7'd073}, '{7'd076, 7'd112, 7'd106, 7'd074}, '{7'd108, 7'd113, 7'd107, 7'd075},
      '{7'd028, 7'd088, 7'd108, 7'd076}, '{7'd060, 7'd089, 7'd109, 7'd077}, '{7'd092, 7'd120, 7'd110, 7'd078}, '{7'd124, 7'd121, 7'd111, 7'd079},
      '{7'd010, 7'd068, 7'd088, 7'd080}, '{7'd042, 7'd069, 7'd089, 7'd081}, '{7'd074, 7'd100, 7'd090, 7'd082}, '{7'd106, 7'd101, 7'd091, 7'd083},
      '{7'd026, 7'd076, 7'd096, 7'd084}, '{7'd058, 7'd077, 7'd097, 7'd085}, '{7'd090, 7'd108, 7'd098, 7'd086}, '{7'd122, 7'd109, 7'd099, 7'd087},
      '{7'd014, 7'd084, 7'd100, 7'd088}, '{7'd046, 7'd085, 7'd101, 7'd089}, '{7'd078, 7'd116, 7'd102, 7'd090}, '{7'd110, 7'd117, 7'd103, 7'd091},
      '{7'd030, 7'd092, 7'd108, 7'd092}, '{7'd062, 7'd093, 7'd109, 7'd093}, '{7'd094, 7'd124, 7'd110, 7'd094}, '{7'd126, 7'd125, 7'd111, 7'd095},
      '{7'd009, 7'd066, 7'd084, 7'd096}, '{7'd041, 7'd067, 7'd085, 7'd097}, '{7'd073, 7'd098, 7'd086, 7'd098}, '{7'd105, 7'd099, 7'd087, 7'd099},
      '{7'd025, 7'd074, 7'd088, 7'd100}, '{7'd057, 7'd075, 7'd089, 7'd101}, '{7'd089, 7'd106, 7'd090, 7'd102}, '{7'd121, 7'd107, 7'd091, 7'd103},
      '{7'd013, 7'd082, 7'd092, 7'd104}, '{7'd045, 7'd083, 7'd093, 7'd105}, '{7'd077, 7'd114, 7'd094, 7'd106}, '{7'd109, 7'd115, 7'd095, 7'd107},
      '{7'd029, 7'd090, 7'd096, 7'd108}, '{7'd061, 7'd091, 7'd097, 7'd109}, '{7'd093, 7'd122, 7'd098, 7'd110}, '{7'd125, 7'd123, 7'd099, 7'd111},
      '{7'd011, 7'd070, 7'd080, 7'd112}, '{7'd043, 7'd071, 7'd081, 7'd113}, '{7'd075, 7'd102, 7'd082, 7'd114}, '{7'd107, 7'd103, 7'd083, 7'd115},
      '{7'd027, 7'd078, 7'd084, 7'd116}, '{7'd059, 7'd079, 7'd085, 7'd117}, '{7'd091, 7'd110, 7'd086, 7'd118}, '{7'd123, 7'd111, 7'd087, 7'd119},
      '{7'd015, 7'd086, 7'd088, 7'd120}, '{7'd047, 7'd087, 7'd089, 7'd121}, '{7'd079, 7'd118, 7'd090, 7'd122}, '{7'd111, 7'd119, 7'd091, 7'd123},
      '{7'd031, 7'd094, 7'd092, 7'd124}, '{7'd063, 7'd095, 7'd093, 7'd125}, '{7'd095, 7'd126, 7'd094, 7'd126}, '{7'd127, 7'd127, 7'd095, 7'd127}
    };

    automatic logic [8-1:0] lut_8lane [0:255][0:3] = '{
      '{8'd000, 8'd000, 8'd000, 8'd000}, '{8'd032, 8'd001, 8'd001, 8'd001}, '{8'd064, 8'd032, 8'd002, 8'd002}, '{8'd096, 8'd033, 8'd003, 8'd003}, '{8'd128, 8'd064, 8'd032, 8'd004}, '{8'd160, 8'd065, 8'd033, 8'd005}, '{8'd192, 8'd096, 8'd034, 8'd006}, '{8'd224, 8'd097, 8'd035, 8'd007},
      '{8'd008, 8'd128, 8'd064, 8'd032}, '{8'd040, 8'd129, 8'd065, 8'd033}, '{8'd072, 8'd160, 8'd066, 8'd034}, '{8'd104, 8'd161, 8'd067, 8'd035}, '{8'd136, 8'd192, 8'd096, 8'd036}, '{8'd168, 8'd193, 8'd097, 8'd037}, '{8'd200, 8'd224, 8'd098, 8'd038}, '{8'd232, 8'd225, 8'd099, 8'd039},
      '{8'd016, 8'd008, 8'd128, 8'd064}, '{8'd048, 8'd009, 8'd129, 8'd065}, '{8'd080, 8'd040, 8'd130, 8'd066}, '{8'd112, 8'd041, 8'd131, 8'd067}, '{8'd144, 8'd072, 8'd160, 8'd068}, '{8'd176, 8'd073, 8'd161, 8'd069}, '{8'd208, 8'd104, 8'd162, 8'd070}, '{8'd240, 8'd105, 8'd163, 8'd071},
      '{8'd024, 8'd136, 8'd192, 8'd096}, '{8'd056, 8'd137, 8'd193, 8'd097}, '{8'd088, 8'd168, 8'd194, 8'd098}, '{8'd120, 8'd169, 8'd195, 8'd099}, '{8'd152, 8'd200, 8'd224, 8'd100}, '{8'd184, 8'd201, 8'd225, 8'd101}, '{8'd216, 8'd232, 8'd226, 8'd102}, '{8'd248, 8'd233, 8'd227, 8'd103},
      '{8'd004, 8'd016, 8'd008, 8'd128}, '{8'd036, 8'd017, 8'd009, 8'd129}, '{8'd068, 8'd048, 8'd010, 8'd130}, '{8'd100, 8'd049, 8'd011, 8'd131}, '{8'd132, 8'd080, 8'd040, 8'd132}, '{8'd164, 8'd081, 8'd041, 8'd133}, '{8'd196, 8'd112, 8'd042, 8'd134}, '{8'd228, 8'd113, 8'd043, 8'd135},
      '{8'd012, 8'd144, 8'd072, 8'd160}, '{8'd044, 8'd145, 8'd073, 8'd161}, '{8'd076, 8'd176, 8'd074, 8'd162}, '{8'd108, 8'd177, 8'd075, 8'd163}, '{8'd140, 8'd208, 8'd104, 8'd164}, '{8'd172, 8'd209, 8'd105, 8'd165}, '{8'd204, 8'd240, 8'd106, 8'd166}, '{8'd236, 8'd241, 8'd107, 8'd167},
      '{8'd020, 8'd024, 8'd136, 8'd192}, '{8'd052, 8'd025, 8'd137, 8'd193}, '{8'd084, 8'd056, 8'd138, 8'd194}, '{8'd116, 8'd057, 8'd139, 8'd195}, '{8'd148, 8'd088, 8'd168, 8'd196}, '{8'd180, 8'd089, 8'd169, 8'd197}, '{8'd212, 8'd120, 8'd170, 8'd198}, '{8'd244, 8'd121, 8'd171, 8'd199},
      '{8'd028, 8'd152, 8'd200, 8'd224}, '{8'd060, 8'd153, 8'd201, 8'd225}, '{8'd092, 8'd184, 8'd202, 8'd226}, '{8'd124, 8'd185, 8'd203, 8'd227}, '{8'd156, 8'd216, 8'd232, 8'd228}, '{8'd188, 8'd217, 8'd233, 8'd229}, '{8'd220, 8'd248, 8'd234, 8'd230}, '{8'd252, 8'd249, 8'd235, 8'd231},
      '{8'd002, 8'd004, 8'd016, 8'd008}, '{8'd034, 8'd005, 8'd017, 8'd009}, '{8'd066, 8'd036, 8'd018, 8'd010}, '{8'd098, 8'd037, 8'd019, 8'd011}, '{8'd130, 8'd068, 8'd048, 8'd012}, '{8'd162, 8'd069, 8'd049, 8'd013}, '{8'd194, 8'd100, 8'd050, 8'd014}, '{8'd226, 8'd101, 8'd051, 8'd015},
      '{8'd010, 8'd132, 8'd080, 8'd040}, '{8'd042, 8'd133, 8'd081, 8'd041}, '{8'd074, 8'd164, 8'd082, 8'd042}, '{8'd106, 8'd165, 8'd083, 8'd043}, '{8'd138, 8'd196, 8'd112, 8'd044}, '{8'd170, 8'd197, 8'd113, 8'd045}, '{8'd202, 8'd228, 8'd114, 8'd046}, '{8'd234, 8'd229, 8'd115, 8'd047},
      '{8'd018, 8'd012, 8'd144, 8'd072}, '{8'd050, 8'd013, 8'd145, 8'd073}, '{8'd082, 8'd044, 8'd146, 8'd074}, '{8'd114, 8'd045, 8'd147, 8'd075}, '{8'd146, 8'd076, 8'd176, 8'd076}, '{8'd178, 8'd077, 8'd177, 8'd077}, '{8'd210, 8'd108, 8'd178, 8'd078}, '{8'd242, 8'd109, 8'd179, 8'd079},
      '{8'd026, 8'd140, 8'd208, 8'd104}, '{8'd058, 8'd141, 8'd209, 8'd105}, '{8'd090, 8'd172, 8'd210, 8'd106}, '{8'd122, 8'd173, 8'd211, 8'd107}, '{8'd154, 8'd204, 8'd240, 8'd108}, '{8'd186, 8'd205, 8'd241, 8'd109}, '{8'd218, 8'd236, 8'd242, 8'd110}, '{8'd250, 8'd237, 8'd243, 8'd111},
      '{8'd006, 8'd020, 8'd024, 8'd136}, '{8'd038, 8'd021, 8'd025, 8'd137}, '{8'd070, 8'd052, 8'd026, 8'd138}, '{8'd102, 8'd053, 8'd027, 8'd139}, '{8'd134, 8'd084, 8'd056, 8'd140}, '{8'd166, 8'd085, 8'd057, 8'd141}, '{8'd198, 8'd116, 8'd058, 8'd142}, '{8'd230, 8'd117, 8'd059, 8'd143},
      '{8'd014, 8'd148, 8'd088, 8'd168}, '{8'd046, 8'd149, 8'd089, 8'd169}, '{8'd078, 8'd180, 8'd090, 8'd170}, '{8'd110, 8'd181, 8'd091, 8'd171}, '{8'd142, 8'd212, 8'd120, 8'd172}, '{8'd174, 8'd213, 8'd121, 8'd173}, '{8'd206, 8'd244, 8'd122, 8'd174}, '{8'd238, 8'd245, 8'd123, 8'd175},
      '{8'd022, 8'd028, 8'd152, 8'd200}, '{8'd054, 8'd029, 8'd153, 8'd201}, '{8'd086, 8'd060, 8'd154, 8'd202}, '{8'd118, 8'd061, 8'd155, 8'd203}, '{8'd150, 8'd092, 8'd184, 8'd204}, '{8'd182, 8'd093, 8'd185, 8'd205}, '{8'd214, 8'd124, 8'd186, 8'd206}, '{8'd246, 8'd125, 8'd187, 8'd207},
      '{8'd030, 8'd156, 8'd216, 8'd232}, '{8'd062, 8'd157, 8'd217, 8'd233}, '{8'd094, 8'd188, 8'd218, 8'd234}, '{8'd126, 8'd189, 8'd219, 8'd235}, '{8'd158, 8'd220, 8'd248, 8'd236}, '{8'd190, 8'd221, 8'd249, 8'd237}, '{8'd222, 8'd252, 8'd250, 8'd238}, '{8'd254, 8'd253, 8'd251, 8'd239},
      '{8'd001, 8'd002, 8'd004, 8'd016}, '{8'd033, 8'd003, 8'd005, 8'd017}, '{8'd065, 8'd034, 8'd006, 8'd018}, '{8'd097, 8'd035, 8'd007, 8'd019}, '{8'd129, 8'd066, 8'd036, 8'd020}, '{8'd161, 8'd067, 8'd037, 8'd021}, '{8'd193, 8'd098, 8'd038, 8'd022}, '{8'd225, 8'd099, 8'd039, 8'd023},
      '{8'd009, 8'd130, 8'd068, 8'd048}, '{8'd041, 8'd131, 8'd069, 8'd049}, '{8'd073, 8'd162, 8'd070, 8'd050}, '{8'd105, 8'd163, 8'd071, 8'd051}, '{8'd137, 8'd194, 8'd100, 8'd052}, '{8'd169, 8'd195, 8'd101, 8'd053}, '{8'd201, 8'd226, 8'd102, 8'd054}, '{8'd233, 8'd227, 8'd103, 8'd055},
      '{8'd017, 8'd010, 8'd132, 8'd080}, '{8'd049, 8'd011, 8'd133, 8'd081}, '{8'd081, 8'd042, 8'd134, 8'd082}, '{8'd113, 8'd043, 8'd135, 8'd083}, '{8'd145, 8'd074, 8'd164, 8'd084}, '{8'd177, 8'd075, 8'd165, 8'd085}, '{8'd209, 8'd106, 8'd166, 8'd086}, '{8'd241, 8'd107, 8'd167, 8'd087},
      '{8'd025, 8'd138, 8'd196, 8'd112}, '{8'd057, 8'd139, 8'd197, 8'd113}, '{8'd089, 8'd170, 8'd198, 8'd114}, '{8'd121, 8'd171, 8'd199, 8'd115}, '{8'd153, 8'd202, 8'd228, 8'd116}, '{8'd185, 8'd203, 8'd229, 8'd117}, '{8'd217, 8'd234, 8'd230, 8'd118}, '{8'd249, 8'd235, 8'd231, 8'd119},
      '{8'd005, 8'd018, 8'd012, 8'd144}, '{8'd037, 8'd019, 8'd013, 8'd145}, '{8'd069, 8'd050, 8'd014, 8'd146}, '{8'd101, 8'd051, 8'd015, 8'd147}, '{8'd133, 8'd082, 8'd044, 8'd148}, '{8'd165, 8'd083, 8'd045, 8'd149}, '{8'd197, 8'd114, 8'd046, 8'd150}, '{8'd229, 8'd115, 8'd047, 8'd151},
      '{8'd013, 8'd146, 8'd076, 8'd176}, '{8'd045, 8'd147, 8'd077, 8'd177}, '{8'd077, 8'd178, 8'd078, 8'd178}, '{8'd109, 8'd179, 8'd079, 8'd179}, '{8'd141, 8'd210, 8'd108, 8'd180}, '{8'd173, 8'd211, 8'd109, 8'd181}, '{8'd205, 8'd242, 8'd110, 8'd182}, '{8'd237, 8'd243, 8'd111, 8'd183},
      '{8'd021, 8'd026, 8'd140, 8'd208}, '{8'd053, 8'd027, 8'd141, 8'd209}, '{8'd085, 8'd058, 8'd142, 8'd210}, '{8'd117, 8'd059, 8'd143, 8'd211}, '{8'd149, 8'd090, 8'd172, 8'd212}, '{8'd181, 8'd091, 8'd173, 8'd213}, '{8'd213, 8'd122, 8'd174, 8'd214}, '{8'd245, 8'd123, 8'd175, 8'd215},
      '{8'd029, 8'd154, 8'd204, 8'd240}, '{8'd061, 8'd155, 8'd205, 8'd241}, '{8'd093, 8'd186, 8'd206, 8'd242}, '{8'd125, 8'd187, 8'd207, 8'd243}, '{8'd157, 8'd218, 8'd236, 8'd244}, '{8'd189, 8'd219, 8'd237, 8'd245}, '{8'd221, 8'd250, 8'd238, 8'd246}, '{8'd253, 8'd251, 8'd239, 8'd247},
      '{8'd003, 8'd006, 8'd020, 8'd024}, '{8'd035, 8'd007, 8'd021, 8'd025}, '{8'd067, 8'd038, 8'd022, 8'd026}, '{8'd099, 8'd039, 8'd023, 8'd027}, '{8'd131, 8'd070, 8'd052, 8'd028}, '{8'd163, 8'd071, 8'd053, 8'd029}, '{8'd195, 8'd102, 8'd054, 8'd030}, '{8'd227, 8'd103, 8'd055, 8'd031},
      '{8'd011, 8'd134, 8'd084, 8'd056}, '{8'd043, 8'd135, 8'd085, 8'd057}, '{8'd075, 8'd166, 8'd086, 8'd058}, '{8'd107, 8'd167, 8'd087, 8'd059}, '{8'd139, 8'd198, 8'd116, 8'd060}, '{8'd171, 8'd199, 8'd117, 8'd061}, '{8'd203, 8'd230, 8'd118, 8'd062}, '{8'd235, 8'd231, 8'd119, 8'd063},
      '{8'd019, 8'd014, 8'd148, 8'd088}, '{8'd051, 8'd015, 8'd149, 8'd089}, '{8'd083, 8'd046, 8'd150, 8'd090}, '{8'd115, 8'd047, 8'd151, 8'd091}, '{8'd147, 8'd078, 8'd180, 8'd092}, '{8'd179, 8'd079, 8'd181, 8'd093}, '{8'd211, 8'd110, 8'd182, 8'd094}, '{8'd243, 8'd111, 8'd183, 8'd095},
      '{8'd027, 8'd142, 8'd212, 8'd120}, '{8'd059, 8'd143, 8'd213, 8'd121}, '{8'd091, 8'd174, 8'd214, 8'd122}, '{8'd123, 8'd175, 8'd215, 8'd123}, '{8'd155, 8'd206, 8'd244, 8'd124}, '{8'd187, 8'd207, 8'd245, 8'd125}, '{8'd219, 8'd238, 8'd246, 8'd126}, '{8'd251, 8'd239, 8'd247, 8'd127},
      '{8'd007, 8'd022, 8'd028, 8'd152}, '{8'd039, 8'd023, 8'd029, 8'd153}, '{8'd071, 8'd054, 8'd030, 8'd154}, '{8'd103, 8'd055, 8'd031, 8'd155}, '{8'd135, 8'd086, 8'd060, 8'd156}, '{8'd167, 8'd087, 8'd061, 8'd157}, '{8'd199, 8'd118, 8'd062, 8'd158}, '{8'd231, 8'd119, 8'd063, 8'd159},
      '{8'd015, 8'd150, 8'd092, 8'd184}, '{8'd047, 8'd151, 8'd093, 8'd185}, '{8'd079, 8'd182, 8'd094, 8'd186}, '{8'd111, 8'd183, 8'd095, 8'd187}, '{8'd143, 8'd214, 8'd124, 8'd188}, '{8'd175, 8'd215, 8'd125, 8'd189}, '{8'd207, 8'd246, 8'd126, 8'd190}, '{8'd239, 8'd247, 8'd127, 8'd191},
      '{8'd023, 8'd030, 8'd156, 8'd216}, '{8'd055, 8'd031, 8'd157, 8'd217}, '{8'd087, 8'd062, 8'd158, 8'd218}, '{8'd119, 8'd063, 8'd159, 8'd219}, '{8'd151, 8'd094, 8'd188, 8'd220}, '{8'd183, 8'd095, 8'd189, 8'd221}, '{8'd215, 8'd126, 8'd190, 8'd222}, '{8'd247, 8'd127, 8'd191, 8'd223},
      '{8'd031, 8'd158, 8'd220, 8'd248}, '{8'd063, 8'd159, 8'd221, 8'd249}, '{8'd095, 8'd190, 8'd222, 8'd250}, '{8'd127, 8'd191, 8'd223, 8'd251}, '{8'd159, 8'd222, 8'd252, 8'd252}, '{8'd191, 8'd223, 8'd253, 8'd253}, '{8'd223, 8'd254, 8'd254, 8'd254}, '{8'd255, 8'd255, 8'd255, 8'd255}
    };

    automatic logic [9-1:0] lut_16lane [0:511][0:3] = '{
      '{9'd000, 9'd000, 9'd000, 9'd000}, '{9'd032, 9'd001, 9'd001, 9'd001}, '{9'd064, 9'd032, 9'd002, 9'd002}, '{9'd096, 9'd033, 9'd003, 9'd003}, '{9'd128, 9'd064, 9'd032, 9'd004}, '{9'd160, 9'd065, 9'd033, 9'd005}, '{9'd192, 9'd096, 9'd034, 9'd006}, '{9'd224, 9'd097, 9'd035, 9'd007},
      '{9'd256, 9'd128, 9'd064, 9'd032}, '{9'd288, 9'd129, 9'd065, 9'd033}, '{9'd320, 9'd160, 9'd066, 9'd034}, '{9'd352, 9'd161, 9'd067, 9'd035}, '{9'd384, 9'd192, 9'd096, 9'd036}, '{9'd416, 9'd193, 9'd097, 9'd037}, '{9'd448, 9'd224, 9'd098, 9'd038}, '{9'd480, 9'd225, 9'd099, 9'd039},
      '{9'd008, 9'd256, 9'd128, 9'd064}, '{9'd040, 9'd257, 9'd129, 9'd065}, '{9'd072, 9'd288, 9'd130, 9'd066}, '{9'd104, 9'd289, 9'd131, 9'd067}, '{9'd136, 9'd320, 9'd160, 9'd068}, '{9'd168, 9'd321, 9'd161, 9'd069}, '{9'd200, 9'd352, 9'd162, 9'd070}, '{9'd232, 9'd353, 9'd163, 9'd071},
      '{9'd264, 9'd384, 9'd192, 9'd096}, '{9'd296, 9'd385, 9'd193, 9'd097}, '{9'd328, 9'd416, 9'd194, 9'd098}, '{9'd360, 9'd417, 9'd195, 9'd099}, '{9'd392, 9'd448, 9'd224, 9'd100}, '{9'd424, 9'd449, 9'd225, 9'd101}, '{9'd456, 9'd480, 9'd226, 9'd102}, '{9'd488, 9'd481, 9'd227, 9'd103},
      '{9'd016, 9'd008, 9'd256, 9'd128}, '{9'd048, 9'd009, 9'd257, 9'd129}, '{9'd080, 9'd040, 9'd258, 9'd130}, '{9'd112, 9'd041, 9'd259, 9'd131}, '{9'd144, 9'd072, 9'd288, 9'd132}, '{9'd176, 9'd073, 9'd289, 9'd133}, '{9'd208, 9'd104, 9'd290, 9'd134}, '{9'd240, 9'd105, 9'd291, 9'd135},
      '{9'd272, 9'd136, 9'd320, 9'd160}, '{9'd304, 9'd137, 9'd321, 9'd161}, '{9'd336, 9'd168, 9'd322, 9'd162}, '{9'd368, 9'd169, 9'd323, 9'd163}, '{9'd400, 9'd200, 9'd352, 9'd164}, '{9'd432, 9'd201, 9'd353, 9'd165}, '{9'd464, 9'd232, 9'd354, 9'd166}, '{9'd496, 9'd233, 9'd355, 9'd167},
      '{9'd024, 9'd264, 9'd384, 9'd192}, '{9'd056, 9'd265, 9'd385, 9'd193}, '{9'd088, 9'd296, 9'd386, 9'd194}, '{9'd120, 9'd297, 9'd387, 9'd195}, '{9'd152, 9'd328, 9'd416, 9'd196}, '{9'd184, 9'd329, 9'd417, 9'd197}, '{9'd216, 9'd360, 9'd418, 9'd198}, '{9'd248, 9'd361, 9'd419, 9'd199},
      '{9'd280, 9'd392, 9'd448, 9'd224}, '{9'd312, 9'd393, 9'd449, 9'd225}, '{9'd344, 9'd424, 9'd450, 9'd226}, '{9'd376, 9'd425, 9'd451, 9'd227}, '{9'd408, 9'd456, 9'd480, 9'd228}, '{9'd440, 9'd457, 9'd481, 9'd229}, '{9'd472, 9'd488, 9'd482, 9'd230}, '{9'd504, 9'd489, 9'd483, 9'd231},
      '{9'd004, 9'd016, 9'd008, 9'd256}, '{9'd036, 9'd017, 9'd009, 9'd257}, '{9'd068, 9'd048, 9'd010, 9'd258}, '{9'd100, 9'd049, 9'd011, 9'd259}, '{9'd132, 9'd080, 9'd040, 9'd260}, '{9'd164, 9'd081, 9'd041, 9'd261}, '{9'd196, 9'd112, 9'd042, 9'd262}, '{9'd228, 9'd113, 9'd043, 9'd263},
      '{9'd260, 9'd144, 9'd072, 9'd288}, '{9'd292, 9'd145, 9'd073, 9'd289}, '{9'd324, 9'd176, 9'd074, 9'd290}, '{9'd356, 9'd177, 9'd075, 9'd291}, '{9'd388, 9'd208, 9'd104, 9'd292}, '{9'd420, 9'd209, 9'd105, 9'd293}, '{9'd452, 9'd240, 9'd106, 9'd294}, '{9'd484, 9'd241, 9'd107, 9'd295},
      '{9'd012, 9'd272, 9'd136, 9'd320}, '{9'd044, 9'd273, 9'd137, 9'd321}, '{9'd076, 9'd304, 9'd138, 9'd322}, '{9'd108, 9'd305, 9'd139, 9'd323}, '{9'd140, 9'd336, 9'd168, 9'd324}, '{9'd172, 9'd337, 9'd169, 9'd325}, '{9'd204, 9'd368, 9'd170, 9'd326}, '{9'd236, 9'd369, 9'd171, 9'd327},
      '{9'd268, 9'd400, 9'd200, 9'd352}, '{9'd300, 9'd401, 9'd201, 9'd353}, '{9'd332, 9'd432, 9'd202, 9'd354}, '{9'd364, 9'd433, 9'd203, 9'd355}, '{9'd396, 9'd464, 9'd232, 9'd356}, '{9'd428, 9'd465, 9'd233, 9'd357}, '{9'd460, 9'd496, 9'd234, 9'd358}, '{9'd492, 9'd497, 9'd235, 9'd359},
      '{9'd020, 9'd024, 9'd264, 9'd384}, '{9'd052, 9'd025, 9'd265, 9'd385}, '{9'd084, 9'd056, 9'd266, 9'd386}, '{9'd116, 9'd057, 9'd267, 9'd387}, '{9'd148, 9'd088, 9'd296, 9'd388}, '{9'd180, 9'd089, 9'd297, 9'd389}, '{9'd212, 9'd120, 9'd298, 9'd390}, '{9'd244, 9'd121, 9'd299, 9'd391},
      '{9'd276, 9'd152, 9'd328, 9'd416}, '{9'd308, 9'd153, 9'd329, 9'd417}, '{9'd340, 9'd184, 9'd330, 9'd418}, '{9'd372, 9'd185, 9'd331, 9'd419}, '{9'd404, 9'd216, 9'd360, 9'd420}, '{9'd436, 9'd217, 9'd361, 9'd421}, '{9'd468, 9'd248, 9'd362, 9'd422}, '{9'd500, 9'd249, 9'd363, 9'd423},
      '{9'd028, 9'd280, 9'd392, 9'd448}, '{9'd060, 9'd281, 9'd393, 9'd449}, '{9'd092, 9'd312, 9'd394, 9'd450}, '{9'd124, 9'd313, 9'd395, 9'd451}, '{9'd156, 9'd344, 9'd424, 9'd452}, '{9'd188, 9'd345, 9'd425, 9'd453}, '{9'd220, 9'd376, 9'd426, 9'd454}, '{9'd252, 9'd377, 9'd427, 9'd455},
      '{9'd284, 9'd408, 9'd456, 9'd480}, '{9'd316, 9'd409, 9'd457, 9'd481}, '{9'd348, 9'd440, 9'd458, 9'd482}, '{9'd380, 9'd441, 9'd459, 9'd483}, '{9'd412, 9'd472, 9'd488, 9'd484}, '{9'd444, 9'd473, 9'd489, 9'd485}, '{9'd476, 9'd504, 9'd490, 9'd486}, '{9'd508, 9'd505, 9'd491, 9'd487},
      '{9'd002, 9'd004, 9'd016, 9'd008}, '{9'd034, 9'd005, 9'd017, 9'd009}, '{9'd066, 9'd036, 9'd018, 9'd010}, '{9'd098, 9'd037, 9'd019, 9'd011}, '{9'd130, 9'd068, 9'd048, 9'd012}, '{9'd162, 9'd069, 9'd049, 9'd013}, '{9'd194, 9'd100, 9'd050, 9'd014}, '{9'd226, 9'd101, 9'd051, 9'd015},
      '{9'd258, 9'd132, 9'd080, 9'd040}, '{9'd290, 9'd133, 9'd081, 9'd041}, '{9'd322, 9'd164, 9'd082, 9'd042}, '{9'd354, 9'd165, 9'd083, 9'd043}, '{9'd386, 9'd196, 9'd112, 9'd044}, '{9'd418, 9'd197, 9'd113, 9'd045}, '{9'd450, 9'd228, 9'd114, 9'd046}, '{9'd482, 9'd229, 9'd115, 9'd047},
      '{9'd010, 9'd260, 9'd144, 9'd072}, '{9'd042, 9'd261, 9'd145, 9'd073}, '{9'd074, 9'd292, 9'd146, 9'd074}, '{9'd106, 9'd293, 9'd147, 9'd075}, '{9'd138, 9'd324, 9'd176, 9'd076}, '{9'd170, 9'd325, 9'd177, 9'd077}, '{9'd202, 9'd356, 9'd178, 9'd078}, '{9'd234, 9'd357, 9'd179, 9'd079},
      '{9'd266, 9'd388, 9'd208, 9'd104}, '{9'd298, 9'd389, 9'd209, 9'd105}, '{9'd330, 9'd420, 9'd210, 9'd106}, '{9'd362, 9'd421, 9'd211, 9'd107}, '{9'd394, 9'd452, 9'd240, 9'd108}, '{9'd426, 9'd453, 9'd241, 9'd109}, '{9'd458, 9'd484, 9'd242, 9'd110}, '{9'd490, 9'd485, 9'd243, 9'd111},
      '{9'd018, 9'd012, 9'd272, 9'd136}, '{9'd050, 9'd013, 9'd273, 9'd137}, '{9'd082, 9'd044, 9'd274, 9'd138}, '{9'd114, 9'd045, 9'd275, 9'd139}, '{9'd146, 9'd076, 9'd304, 9'd140}, '{9'd178, 9'd077, 9'd305, 9'd141}, '{9'd210, 9'd108, 9'd306, 9'd142}, '{9'd242, 9'd109, 9'd307, 9'd143},
      '{9'd274, 9'd140, 9'd336, 9'd168}, '{9'd306, 9'd141, 9'd337, 9'd169}, '{9'd338, 9'd172, 9'd338, 9'd170}, '{9'd370, 9'd173, 9'd339, 9'd171}, '{9'd402, 9'd204, 9'd368, 9'd172}, '{9'd434, 9'd205, 9'd369, 9'd173}, '{9'd466, 9'd236, 9'd370, 9'd174}, '{9'd498, 9'd237, 9'd371, 9'd175},
      '{9'd026, 9'd268, 9'd400, 9'd200}, '{9'd058, 9'd269, 9'd401, 9'd201}, '{9'd090, 9'd300, 9'd402, 9'd202}, '{9'd122, 9'd301, 9'd403, 9'd203}, '{9'd154, 9'd332, 9'd432, 9'd204}, '{9'd186, 9'd333, 9'd433, 9'd205}, '{9'd218, 9'd364, 9'd434, 9'd206}, '{9'd250, 9'd365, 9'd435, 9'd207},
      '{9'd282, 9'd396, 9'd464, 9'd232}, '{9'd314, 9'd397, 9'd465, 9'd233}, '{9'd346, 9'd428, 9'd466, 9'd234}, '{9'd378, 9'd429, 9'd467, 9'd235}, '{9'd410, 9'd460, 9'd496, 9'd236}, '{9'd442, 9'd461, 9'd497, 9'd237}, '{9'd474, 9'd492, 9'd498, 9'd238}, '{9'd506, 9'd493, 9'd499, 9'd239},
      '{9'd006, 9'd020, 9'd024, 9'd264}, '{9'd038, 9'd021, 9'd025, 9'd265}, '{9'd070, 9'd052, 9'd026, 9'd266}, '{9'd102, 9'd053, 9'd027, 9'd267}, '{9'd134, 9'd084, 9'd056, 9'd268}, '{9'd166, 9'd085, 9'd057, 9'd269}, '{9'd198, 9'd116, 9'd058, 9'd270}, '{9'd230, 9'd117, 9'd059, 9'd271},
      '{9'd262, 9'd148, 9'd088, 9'd296}, '{9'd294, 9'd149, 9'd089, 9'd297}, '{9'd326, 9'd180, 9'd090, 9'd298}, '{9'd358, 9'd181, 9'd091, 9'd299}, '{9'd390, 9'd212, 9'd120, 9'd300}, '{9'd422, 9'd213, 9'd121, 9'd301}, '{9'd454, 9'd244, 9'd122, 9'd302}, '{9'd486, 9'd245, 9'd123, 9'd303},
      '{9'd014, 9'd276, 9'd152, 9'd328}, '{9'd046, 9'd277, 9'd153, 9'd329}, '{9'd078, 9'd308, 9'd154, 9'd330}, '{9'd110, 9'd309, 9'd155, 9'd331}, '{9'd142, 9'd340, 9'd184, 9'd332}, '{9'd174, 9'd341, 9'd185, 9'd333}, '{9'd206, 9'd372, 9'd186, 9'd334}, '{9'd238, 9'd373, 9'd187, 9'd335},
      '{9'd270, 9'd404, 9'd216, 9'd360}, '{9'd302, 9'd405, 9'd217, 9'd361}, '{9'd334, 9'd436, 9'd218, 9'd362}, '{9'd366, 9'd437, 9'd219, 9'd363}, '{9'd398, 9'd468, 9'd248, 9'd364}, '{9'd430, 9'd469, 9'd249, 9'd365}, '{9'd462, 9'd500, 9'd250, 9'd366}, '{9'd494, 9'd501, 9'd251, 9'd367},
      '{9'd022, 9'd028, 9'd280, 9'd392}, '{9'd054, 9'd029, 9'd281, 9'd393}, '{9'd086, 9'd060, 9'd282, 9'd394}, '{9'd118, 9'd061, 9'd283, 9'd395}, '{9'd150, 9'd092, 9'd312, 9'd396}, '{9'd182, 9'd093, 9'd313, 9'd397}, '{9'd214, 9'd124, 9'd314, 9'd398}, '{9'd246, 9'd125, 9'd315, 9'd399},
      '{9'd278, 9'd156, 9'd344, 9'd424}, '{9'd310, 9'd157, 9'd345, 9'd425}, '{9'd342, 9'd188, 9'd346, 9'd426}, '{9'd374, 9'd189, 9'd347, 9'd427}, '{9'd406, 9'd220, 9'd376, 9'd428}, '{9'd438, 9'd221, 9'd377, 9'd429}, '{9'd470, 9'd252, 9'd378, 9'd430}, '{9'd502, 9'd253, 9'd379, 9'd431},
      '{9'd030, 9'd284, 9'd408, 9'd456}, '{9'd062, 9'd285, 9'd409, 9'd457}, '{9'd094, 9'd316, 9'd410, 9'd458}, '{9'd126, 9'd317, 9'd411, 9'd459}, '{9'd158, 9'd348, 9'd440, 9'd460}, '{9'd190, 9'd349, 9'd441, 9'd461}, '{9'd222, 9'd380, 9'd442, 9'd462}, '{9'd254, 9'd381, 9'd443, 9'd463},
      '{9'd286, 9'd412, 9'd472, 9'd488}, '{9'd318, 9'd413, 9'd473, 9'd489}, '{9'd350, 9'd444, 9'd474, 9'd490}, '{9'd382, 9'd445, 9'd475, 9'd491}, '{9'd414, 9'd476, 9'd504, 9'd492}, '{9'd446, 9'd477, 9'd505, 9'd493}, '{9'd478, 9'd508, 9'd506, 9'd494}, '{9'd510, 9'd509, 9'd507, 9'd495},
      '{9'd001, 9'd002, 9'd004, 9'd016}, '{9'd033, 9'd003, 9'd005, 9'd017}, '{9'd065, 9'd034, 9'd006, 9'd018}, '{9'd097, 9'd035, 9'd007, 9'd019}, '{9'd129, 9'd066, 9'd036, 9'd020}, '{9'd161, 9'd067, 9'd037, 9'd021}, '{9'd193, 9'd098, 9'd038, 9'd022}, '{9'd225, 9'd099, 9'd039, 9'd023},
      '{9'd257, 9'd130, 9'd068, 9'd048}, '{9'd289, 9'd131, 9'd069, 9'd049}, '{9'd321, 9'd162, 9'd070, 9'd050}, '{9'd353, 9'd163, 9'd071, 9'd051}, '{9'd385, 9'd194, 9'd100, 9'd052}, '{9'd417, 9'd195, 9'd101, 9'd053}, '{9'd449, 9'd226, 9'd102, 9'd054}, '{9'd481, 9'd227, 9'd103, 9'd055},
      '{9'd009, 9'd258, 9'd132, 9'd080}, '{9'd041, 9'd259, 9'd133, 9'd081}, '{9'd073, 9'd290, 9'd134, 9'd082}, '{9'd105, 9'd291, 9'd135, 9'd083}, '{9'd137, 9'd322, 9'd164, 9'd084}, '{9'd169, 9'd323, 9'd165, 9'd085}, '{9'd201, 9'd354, 9'd166, 9'd086}, '{9'd233, 9'd355, 9'd167, 9'd087},
      '{9'd265, 9'd386, 9'd196, 9'd112}, '{9'd297, 9'd387, 9'd197, 9'd113}, '{9'd329, 9'd418, 9'd198, 9'd114}, '{9'd361, 9'd419, 9'd199, 9'd115}, '{9'd393, 9'd450, 9'd228, 9'd116}, '{9'd425, 9'd451, 9'd229, 9'd117}, '{9'd457, 9'd482, 9'd230, 9'd118}, '{9'd489, 9'd483, 9'd231, 9'd119},
      '{9'd017, 9'd010, 9'd260, 9'd144}, '{9'd049, 9'd011, 9'd261, 9'd145}, '{9'd081, 9'd042, 9'd262, 9'd146}, '{9'd113, 9'd043, 9'd263, 9'd147}, '{9'd145, 9'd074, 9'd292, 9'd148}, '{9'd177, 9'd075, 9'd293, 9'd149}, '{9'd209, 9'd106, 9'd294, 9'd150}, '{9'd241, 9'd107, 9'd295, 9'd151},
      '{9'd273, 9'd138, 9'd324, 9'd176}, '{9'd305, 9'd139, 9'd325, 9'd177}, '{9'd337, 9'd170, 9'd326, 9'd178}, '{9'd369, 9'd171, 9'd327, 9'd179}, '{9'd401, 9'd202, 9'd356, 9'd180}, '{9'd433, 9'd203, 9'd357, 9'd181}, '{9'd465, 9'd234, 9'd358, 9'd182}, '{9'd497, 9'd235, 9'd359, 9'd183},
      '{9'd025, 9'd266, 9'd388, 9'd208}, '{9'd057, 9'd267, 9'd389, 9'd209}, '{9'd089, 9'd298, 9'd390, 9'd210}, '{9'd121, 9'd299, 9'd391, 9'd211}, '{9'd153, 9'd330, 9'd420, 9'd212}, '{9'd185, 9'd331, 9'd421, 9'd213}, '{9'd217, 9'd362, 9'd422, 9'd214}, '{9'd249, 9'd363, 9'd423, 9'd215},
      '{9'd281, 9'd394, 9'd452, 9'd240}, '{9'd313, 9'd395, 9'd453, 9'd241}, '{9'd345, 9'd426, 9'd454, 9'd242}, '{9'd377, 9'd427, 9'd455, 9'd243}, '{9'd409, 9'd458, 9'd484, 9'd244}, '{9'd441, 9'd459, 9'd485, 9'd245}, '{9'd473, 9'd490, 9'd486, 9'd246}, '{9'd505, 9'd491, 9'd487, 9'd247},
      '{9'd005, 9'd018, 9'd012, 9'd272}, '{9'd037, 9'd019, 9'd013, 9'd273}, '{9'd069, 9'd050, 9'd014, 9'd274}, '{9'd101, 9'd051, 9'd015, 9'd275}, '{9'd133, 9'd082, 9'd044, 9'd276}, '{9'd165, 9'd083, 9'd045, 9'd277}, '{9'd197, 9'd114, 9'd046, 9'd278}, '{9'd229, 9'd115, 9'd047, 9'd279},
      '{9'd261, 9'd146, 9'd076, 9'd304}, '{9'd293, 9'd147, 9'd077, 9'd305}, '{9'd325, 9'd178, 9'd078, 9'd306}, '{9'd357, 9'd179, 9'd079, 9'd307}, '{9'd389, 9'd210, 9'd108, 9'd308}, '{9'd421, 9'd211, 9'd109, 9'd309}, '{9'd453, 9'd242, 9'd110, 9'd310}, '{9'd485, 9'd243, 9'd111, 9'd311},
      '{9'd013, 9'd274, 9'd140, 9'd336}, '{9'd045, 9'd275, 9'd141, 9'd337}, '{9'd077, 9'd306, 9'd142, 9'd338}, '{9'd109, 9'd307, 9'd143, 9'd339}, '{9'd141, 9'd338, 9'd172, 9'd340}, '{9'd173, 9'd339, 9'd173, 9'd341}, '{9'd205, 9'd370, 9'd174, 9'd342}, '{9'd237, 9'd371, 9'd175, 9'd343},
      '{9'd269, 9'd402, 9'd204, 9'd368}, '{9'd301, 9'd403, 9'd205, 9'd369}, '{9'd333, 9'd434, 9'd206, 9'd370}, '{9'd365, 9'd435, 9'd207, 9'd371}, '{9'd397, 9'd466, 9'd236, 9'd372}, '{9'd429, 9'd467, 9'd237, 9'd373}, '{9'd461, 9'd498, 9'd238, 9'd374}, '{9'd493, 9'd499, 9'd239, 9'd375},
      '{9'd021, 9'd026, 9'd268, 9'd400}, '{9'd053, 9'd027, 9'd269, 9'd401}, '{9'd085, 9'd058, 9'd270, 9'd402}, '{9'd117, 9'd059, 9'd271, 9'd403}, '{9'd149, 9'd090, 9'd300, 9'd404}, '{9'd181, 9'd091, 9'd301, 9'd405}, '{9'd213, 9'd122, 9'd302, 9'd406}, '{9'd245, 9'd123, 9'd303, 9'd407},
      '{9'd277, 9'd154, 9'd332, 9'd432}, '{9'd309, 9'd155, 9'd333, 9'd433}, '{9'd341, 9'd186, 9'd334, 9'd434}, '{9'd373, 9'd187, 9'd335, 9'd435}, '{9'd405, 9'd218, 9'd364, 9'd436}, '{9'd437, 9'd219, 9'd365, 9'd437}, '{9'd469, 9'd250, 9'd366, 9'd438}, '{9'd501, 9'd251, 9'd367, 9'd439},
      '{9'd029, 9'd282, 9'd396, 9'd464}, '{9'd061, 9'd283, 9'd397, 9'd465}, '{9'd093, 9'd314, 9'd398, 9'd466}, '{9'd125, 9'd315, 9'd399, 9'd467}, '{9'd157, 9'd346, 9'd428, 9'd468}, '{9'd189, 9'd347, 9'd429, 9'd469}, '{9'd221, 9'd378, 9'd430, 9'd470}, '{9'd253, 9'd379, 9'd431, 9'd471},
      '{9'd285, 9'd410, 9'd460, 9'd496}, '{9'd317, 9'd411, 9'd461, 9'd497}, '{9'd349, 9'd442, 9'd462, 9'd498}, '{9'd381, 9'd443, 9'd463, 9'd499}, '{9'd413, 9'd474, 9'd492, 9'd500}, '{9'd445, 9'd475, 9'd493, 9'd501}, '{9'd477, 9'd506, 9'd494, 9'd502}, '{9'd509, 9'd507, 9'd495, 9'd503},
      '{9'd003, 9'd006, 9'd020, 9'd024}, '{9'd035, 9'd007, 9'd021, 9'd025}, '{9'd067, 9'd038, 9'd022, 9'd026}, '{9'd099, 9'd039, 9'd023, 9'd027}, '{9'd131, 9'd070, 9'd052, 9'd028}, '{9'd163, 9'd071, 9'd053, 9'd029}, '{9'd195, 9'd102, 9'd054, 9'd030}, '{9'd227, 9'd103, 9'd055, 9'd031},
      '{9'd259, 9'd134, 9'd084, 9'd056}, '{9'd291, 9'd135, 9'd085, 9'd057}, '{9'd323, 9'd166, 9'd086, 9'd058}, '{9'd355, 9'd167, 9'd087, 9'd059}, '{9'd387, 9'd198, 9'd116, 9'd060}, '{9'd419, 9'd199, 9'd117, 9'd061}, '{9'd451, 9'd230, 9'd118, 9'd062}, '{9'd483, 9'd231, 9'd119, 9'd063},
      '{9'd011, 9'd262, 9'd148, 9'd088}, '{9'd043, 9'd263, 9'd149, 9'd089}, '{9'd075, 9'd294, 9'd150, 9'd090}, '{9'd107, 9'd295, 9'd151, 9'd091}, '{9'd139, 9'd326, 9'd180, 9'd092}, '{9'd171, 9'd327, 9'd181, 9'd093}, '{9'd203, 9'd358, 9'd182, 9'd094}, '{9'd235, 9'd359, 9'd183, 9'd095},
      '{9'd267, 9'd390, 9'd212, 9'd120}, '{9'd299, 9'd391, 9'd213, 9'd121}, '{9'd331, 9'd422, 9'd214, 9'd122}, '{9'd363, 9'd423, 9'd215, 9'd123}, '{9'd395, 9'd454, 9'd244, 9'd124}, '{9'd427, 9'd455, 9'd245, 9'd125}, '{9'd459, 9'd486, 9'd246, 9'd126}, '{9'd491, 9'd487, 9'd247, 9'd127},
      '{9'd019, 9'd014, 9'd276, 9'd152}, '{9'd051, 9'd015, 9'd277, 9'd153}, '{9'd083, 9'd046, 9'd278, 9'd154}, '{9'd115, 9'd047, 9'd279, 9'd155}, '{9'd147, 9'd078, 9'd308, 9'd156}, '{9'd179, 9'd079, 9'd309, 9'd157}, '{9'd211, 9'd110, 9'd310, 9'd158}, '{9'd243, 9'd111, 9'd311, 9'd159},
      '{9'd275, 9'd142, 9'd340, 9'd184}, '{9'd307, 9'd143, 9'd341, 9'd185}, '{9'd339, 9'd174, 9'd342, 9'd186}, '{9'd371, 9'd175, 9'd343, 9'd187}, '{9'd403, 9'd206, 9'd372, 9'd188}, '{9'd435, 9'd207, 9'd373, 9'd189}, '{9'd467, 9'd238, 9'd374, 9'd190}, '{9'd499, 9'd239, 9'd375, 9'd191},
      '{9'd027, 9'd270, 9'd404, 9'd216}, '{9'd059, 9'd271, 9'd405, 9'd217}, '{9'd091, 9'd302, 9'd406, 9'd218}, '{9'd123, 9'd303, 9'd407, 9'd219}, '{9'd155, 9'd334, 9'd436, 9'd220}, '{9'd187, 9'd335, 9'd437, 9'd221}, '{9'd219, 9'd366, 9'd438, 9'd222}, '{9'd251, 9'd367, 9'd439, 9'd223},
      '{9'd283, 9'd398, 9'd468, 9'd248}, '{9'd315, 9'd399, 9'd469, 9'd249}, '{9'd347, 9'd430, 9'd470, 9'd250}, '{9'd379, 9'd431, 9'd471, 9'd251}, '{9'd411, 9'd462, 9'd500, 9'd252}, '{9'd443, 9'd463, 9'd501, 9'd253}, '{9'd475, 9'd494, 9'd502, 9'd254}, '{9'd507, 9'd495, 9'd503, 9'd255},
      '{9'd007, 9'd022, 9'd028, 9'd280}, '{9'd039, 9'd023, 9'd029, 9'd281}, '{9'd071, 9'd054, 9'd030, 9'd282}, '{9'd103, 9'd055, 9'd031, 9'd283}, '{9'd135, 9'd086, 9'd060, 9'd284}, '{9'd167, 9'd087, 9'd061, 9'd285}, '{9'd199, 9'd118, 9'd062, 9'd286}, '{9'd231, 9'd119, 9'd063, 9'd287},
      '{9'd263, 9'd150, 9'd092, 9'd312}, '{9'd295, 9'd151, 9'd093, 9'd313}, '{9'd327, 9'd182, 9'd094, 9'd314}, '{9'd359, 9'd183, 9'd095, 9'd315}, '{9'd391, 9'd214, 9'd124, 9'd316}, '{9'd423, 9'd215, 9'd125, 9'd317}, '{9'd455, 9'd246, 9'd126, 9'd318}, '{9'd487, 9'd247, 9'd127, 9'd319},
      '{9'd015, 9'd278, 9'd156, 9'd344}, '{9'd047, 9'd279, 9'd157, 9'd345}, '{9'd079, 9'd310, 9'd158, 9'd346}, '{9'd111, 9'd311, 9'd159, 9'd347}, '{9'd143, 9'd342, 9'd188, 9'd348}, '{9'd175, 9'd343, 9'd189, 9'd349}, '{9'd207, 9'd374, 9'd190, 9'd350}, '{9'd239, 9'd375, 9'd191, 9'd351},
      '{9'd271, 9'd406, 9'd220, 9'd376}, '{9'd303, 9'd407, 9'd221, 9'd377}, '{9'd335, 9'd438, 9'd222, 9'd378}, '{9'd367, 9'd439, 9'd223, 9'd379}, '{9'd399, 9'd470, 9'd252, 9'd380}, '{9'd431, 9'd471, 9'd253, 9'd381}, '{9'd463, 9'd502, 9'd254, 9'd382}, '{9'd495, 9'd503, 9'd255, 9'd383},
      '{9'd023, 9'd030, 9'd284, 9'd408}, '{9'd055, 9'd031, 9'd285, 9'd409}, '{9'd087, 9'd062, 9'd286, 9'd410}, '{9'd119, 9'd063, 9'd287, 9'd411}, '{9'd151, 9'd094, 9'd316, 9'd412}, '{9'd183, 9'd095, 9'd317, 9'd413}, '{9'd215, 9'd126, 9'd318, 9'd414}, '{9'd247, 9'd127, 9'd319, 9'd415},
      '{9'd279, 9'd158, 9'd348, 9'd440}, '{9'd311, 9'd159, 9'd349, 9'd441}, '{9'd343, 9'd190, 9'd350, 9'd442}, '{9'd375, 9'd191, 9'd351, 9'd443}, '{9'd407, 9'd222, 9'd380, 9'd444}, '{9'd439, 9'd223, 9'd381, 9'd445}, '{9'd471, 9'd254, 9'd382, 9'd446}, '{9'd503, 9'd255, 9'd383, 9'd447},
      '{9'd031, 9'd286, 9'd412, 9'd472}, '{9'd063, 9'd287, 9'd413, 9'd473}, '{9'd095, 9'd318, 9'd414, 9'd474}, '{9'd127, 9'd319, 9'd415, 9'd475}, '{9'd159, 9'd350, 9'd444, 9'd476}, '{9'd191, 9'd351, 9'd445, 9'd477}, '{9'd223, 9'd382, 9'd446, 9'd478}, '{9'd255, 9'd383, 9'd447, 9'd479},
      '{9'd287, 9'd414, 9'd476, 9'd504}, '{9'd319, 9'd415, 9'd477, 9'd505}, '{9'd351, 9'd446, 9'd478, 9'd506}, '{9'd383, 9'd447, 9'd479, 9'd507}, '{9'd415, 9'd478, 9'd508, 9'd508}, '{9'd447, 9'd479, 9'd509, 9'd509}, '{9'd479, 9'd510, 9'd510, 9'd510}, '{9'd511, 9'd511, 9'd511, 9'd511}
    };

	unique case (NrLanes)
      1 : return lut_1lane [seqNbIdx][ew];
      2 : return lut_2lane [seqNbIdx][ew];
      4 : return lut_4lane [seqNbIdx][ew];
      8 : return lut_8lane [seqNbIdx][ew];
      16: return lut_16lane[seqNbIdx][ew];
      default: return 0;
	  endcase
  endfunction

  function automatic logic [{$clog2(riva_pkg::DLEN*riva_pkg::MaxNrLanes/4)}-1:0] query_shf_idx_2d_cln(input int NrLanes, input int seqNbIdx, input riscv_mv_pkg::vew_e ew);
    automatic logic [5-1:0] lut_1lane [0:31][0:3] = '{
      '{5'd000, 5'd000, 5'd000, 5'd000}, '{5'd008, 5'd001, 5'd001, 5'd001}, '{5'd016, 5'd008, 5'd002, 5'd002}, '{5'd024, 5'd009, 5'd003, 5'd003}, '{5'd004, 5'd016, 5'd008, 5'd004}, '{5'd012, 5'd017, 5'd009, 5'd005}, '{5'd020, 5'd024, 5'd010, 5'd006}, '{5'd028, 5'd025, 5'd011, 5'd007},
      '{5'd002, 5'd004, 5'd016, 5'd008}, '{5'd010, 5'd005, 5'd017, 5'd009}, '{5'd018, 5'd012, 5'd018, 5'd010}, '{5'd026, 5'd013, 5'd019, 5'd011}, '{5'd006, 5'd020, 5'd024, 5'd012}, '{5'd014, 5'd021, 5'd025, 5'd013}, '{5'd022, 5'd028, 5'd026, 5'd014}, '{5'd030, 5'd029, 5'd027, 5'd015},
      '{5'd001, 5'd002, 5'd004, 5'd016}, '{5'd009, 5'd003, 5'd005, 5'd017}, '{5'd017, 5'd010, 5'd006, 5'd018}, '{5'd025, 5'd011, 5'd007, 5'd019}, '{5'd005, 5'd018, 5'd012, 5'd020}, '{5'd013, 5'd019, 5'd013, 5'd021}, '{5'd021, 5'd026, 5'd014, 5'd022}, '{5'd029, 5'd027, 5'd015, 5'd023},
      '{5'd003, 5'd006, 5'd020, 5'd024}, '{5'd011, 5'd007, 5'd021, 5'd025}, '{5'd019, 5'd014, 5'd022, 5'd026}, '{5'd027, 5'd015, 5'd023, 5'd027}, '{5'd007, 5'd022, 5'd028, 5'd028}, '{5'd015, 5'd023, 5'd029, 5'd029}, '{5'd023, 5'd030, 5'd030, 5'd030}, '{5'd031, 5'd031, 5'd031, 5'd031}
    };

    automatic logic [6-1:0] lut_2lane [0:63][0:3] = '{
      '{6'd000, 6'd000, 6'd000, 6'd000}, '{6'd008, 6'd001, 6'd001, 6'd001}, '{6'd016, 6'd008, 6'd002, 6'd002}, '{6'd024, 6'd009, 6'd003, 6'd003}, '{6'd004, 6'd016, 6'd008, 6'd004}, '{6'd012, 6'd017, 6'd009, 6'd005}, '{6'd020, 6'd024, 6'd010, 6'd006}, '{6'd028, 6'd025, 6'd011, 6'd007},
      '{6'd002, 6'd004, 6'd016, 6'd008}, '{6'd010, 6'd005, 6'd017, 6'd009}, '{6'd018, 6'd012, 6'd018, 6'd010}, '{6'd026, 6'd013, 6'd019, 6'd011}, '{6'd006, 6'd020, 6'd024, 6'd012}, '{6'd014, 6'd021, 6'd025, 6'd013}, '{6'd022, 6'd028, 6'd026, 6'd014}, '{6'd030, 6'd029, 6'd027, 6'd015},
      '{6'd001, 6'd002, 6'd004, 6'd016}, '{6'd009, 6'd003, 6'd005, 6'd017}, '{6'd017, 6'd010, 6'd006, 6'd018}, '{6'd025, 6'd011, 6'd007, 6'd019}, '{6'd005, 6'd018, 6'd012, 6'd020}, '{6'd013, 6'd019, 6'd013, 6'd021}, '{6'd021, 6'd026, 6'd014, 6'd022}, '{6'd029, 6'd027, 6'd015, 6'd023},
      '{6'd003, 6'd006, 6'd020, 6'd024}, '{6'd011, 6'd007, 6'd021, 6'd025}, '{6'd019, 6'd014, 6'd022, 6'd026}, '{6'd027, 6'd015, 6'd023, 6'd027}, '{6'd007, 6'd022, 6'd028, 6'd028}, '{6'd015, 6'd023, 6'd029, 6'd029}, '{6'd023, 6'd030, 6'd030, 6'd030}, '{6'd031, 6'd031, 6'd031, 6'd031},
      '{6'd032, 6'd032, 6'd032, 6'd032}, '{6'd040, 6'd033, 6'd033, 6'd033}, '{6'd048, 6'd040, 6'd034, 6'd034}, '{6'd056, 6'd041, 6'd035, 6'd035}, '{6'd036, 6'd048, 6'd040, 6'd036}, '{6'd044, 6'd049, 6'd041, 6'd037}, '{6'd052, 6'd056, 6'd042, 6'd038}, '{6'd060, 6'd057, 6'd043, 6'd039},
      '{6'd034, 6'd036, 6'd048, 6'd040}, '{6'd042, 6'd037, 6'd049, 6'd041}, '{6'd050, 6'd044, 6'd050, 6'd042}, '{6'd058, 6'd045, 6'd051, 6'd043}, '{6'd038, 6'd052, 6'd056, 6'd044}, '{6'd046, 6'd053, 6'd057, 6'd045}, '{6'd054, 6'd060, 6'd058, 6'd046}, '{6'd062, 6'd061, 6'd059, 6'd047},
      '{6'd033, 6'd034, 6'd036, 6'd048}, '{6'd041, 6'd035, 6'd037, 6'd049}, '{6'd049, 6'd042, 6'd038, 6'd050}, '{6'd057, 6'd043, 6'd039, 6'd051}, '{6'd037, 6'd050, 6'd044, 6'd052}, '{6'd045, 6'd051, 6'd045, 6'd053}, '{6'd053, 6'd058, 6'd046, 6'd054}, '{6'd061, 6'd059, 6'd047, 6'd055},
      '{6'd035, 6'd038, 6'd052, 6'd056}, '{6'd043, 6'd039, 6'd053, 6'd057}, '{6'd051, 6'd046, 6'd054, 6'd058}, '{6'd059, 6'd047, 6'd055, 6'd059}, '{6'd039, 6'd054, 6'd060, 6'd060}, '{6'd047, 6'd055, 6'd061, 6'd061}, '{6'd055, 6'd062, 6'd062, 6'd062}, '{6'd063, 6'd063, 6'd063, 6'd063}
    };

    automatic logic [7-1:0] lut_4lane [0:127][0:3] = '{
      '{7'd000, 7'd000, 7'd000, 7'd000}, '{7'd008, 7'd001, 7'd001, 7'd001}, '{7'd016, 7'd008, 7'd002, 7'd002}, '{7'd024, 7'd009, 7'd003, 7'd003}, '{7'd004, 7'd016, 7'd008, 7'd004}, '{7'd012, 7'd017, 7'd009, 7'd005}, '{7'd020, 7'd024, 7'd010, 7'd006}, '{7'd028, 7'd025, 7'd011, 7'd007},
      '{7'd002, 7'd004, 7'd016, 7'd008}, '{7'd010, 7'd005, 7'd017, 7'd009}, '{7'd018, 7'd012, 7'd018, 7'd010}, '{7'd026, 7'd013, 7'd019, 7'd011}, '{7'd006, 7'd020, 7'd024, 7'd012}, '{7'd014, 7'd021, 7'd025, 7'd013}, '{7'd022, 7'd028, 7'd026, 7'd014}, '{7'd030, 7'd029, 7'd027, 7'd015},
      '{7'd001, 7'd002, 7'd004, 7'd016}, '{7'd009, 7'd003, 7'd005, 7'd017}, '{7'd017, 7'd010, 7'd006, 7'd018}, '{7'd025, 7'd011, 7'd007, 7'd019}, '{7'd005, 7'd018, 7'd012, 7'd020}, '{7'd013, 7'd019, 7'd013, 7'd021}, '{7'd021, 7'd026, 7'd014, 7'd022}, '{7'd029, 7'd027, 7'd015, 7'd023},
      '{7'd003, 7'd006, 7'd020, 7'd024}, '{7'd011, 7'd007, 7'd021, 7'd025}, '{7'd019, 7'd014, 7'd022, 7'd026}, '{7'd027, 7'd015, 7'd023, 7'd027}, '{7'd007, 7'd022, 7'd028, 7'd028}, '{7'd015, 7'd023, 7'd029, 7'd029}, '{7'd023, 7'd030, 7'd030, 7'd030}, '{7'd031, 7'd031, 7'd031, 7'd031},
      '{7'd032, 7'd032, 7'd032, 7'd032}, '{7'd040, 7'd033, 7'd033, 7'd033}, '{7'd048, 7'd040, 7'd034, 7'd034}, '{7'd056, 7'd041, 7'd035, 7'd035}, '{7'd036, 7'd048, 7'd040, 7'd036}, '{7'd044, 7'd049, 7'd041, 7'd037}, '{7'd052, 7'd056, 7'd042, 7'd038}, '{7'd060, 7'd057, 7'd043, 7'd039},
      '{7'd034, 7'd036, 7'd048, 7'd040}, '{7'd042, 7'd037, 7'd049, 7'd041}, '{7'd050, 7'd044, 7'd050, 7'd042}, '{7'd058, 7'd045, 7'd051, 7'd043}, '{7'd038, 7'd052, 7'd056, 7'd044}, '{7'd046, 7'd053, 7'd057, 7'd045}, '{7'd054, 7'd060, 7'd058, 7'd046}, '{7'd062, 7'd061, 7'd059, 7'd047},
      '{7'd033, 7'd034, 7'd036, 7'd048}, '{7'd041, 7'd035, 7'd037, 7'd049}, '{7'd049, 7'd042, 7'd038, 7'd050}, '{7'd057, 7'd043, 7'd039, 7'd051}, '{7'd037, 7'd050, 7'd044, 7'd052}, '{7'd045, 7'd051, 7'd045, 7'd053}, '{7'd053, 7'd058, 7'd046, 7'd054}, '{7'd061, 7'd059, 7'd047, 7'd055},
      '{7'd035, 7'd038, 7'd052, 7'd056}, '{7'd043, 7'd039, 7'd053, 7'd057}, '{7'd051, 7'd046, 7'd054, 7'd058}, '{7'd059, 7'd047, 7'd055, 7'd059}, '{7'd039, 7'd054, 7'd060, 7'd060}, '{7'd047, 7'd055, 7'd061, 7'd061}, '{7'd055, 7'd062, 7'd062, 7'd062}, '{7'd063, 7'd063, 7'd063, 7'd063},
      '{7'd064, 7'd064, 7'd064, 7'd064}, '{7'd072, 7'd065, 7'd065, 7'd065}, '{7'd080, 7'd072, 7'd066, 7'd066}, '{7'd088, 7'd073, 7'd067, 7'd067}, '{7'd068, 7'd080, 7'd072, 7'd068}, '{7'd076, 7'd081, 7'd073, 7'd069}, '{7'd084, 7'd088, 7'd074, 7'd070}, '{7'd092, 7'd089, 7'd075, 7'd071},
      '{7'd066, 7'd068, 7'd080, 7'd072}, '{7'd074, 7'd069, 7'd081, 7'd073}, '{7'd082, 7'd076, 7'd082, 7'd074}, '{7'd090, 7'd077, 7'd083, 7'd075}, '{7'd070, 7'd084, 7'd088, 7'd076}, '{7'd078, 7'd085, 7'd089, 7'd077}, '{7'd086, 7'd092, 7'd090, 7'd078}, '{7'd094, 7'd093, 7'd091, 7'd079},
      '{7'd065, 7'd066, 7'd068, 7'd080}, '{7'd073, 7'd067, 7'd069, 7'd081}, '{7'd081, 7'd074, 7'd070, 7'd082}, '{7'd089, 7'd075, 7'd071, 7'd083}, '{7'd069, 7'd082, 7'd076, 7'd084}, '{7'd077, 7'd083, 7'd077, 7'd085}, '{7'd085, 7'd090, 7'd078, 7'd086}, '{7'd093, 7'd091, 7'd079, 7'd087},
      '{7'd067, 7'd070, 7'd084, 7'd088}, '{7'd075, 7'd071, 7'd085, 7'd089}, '{7'd083, 7'd078, 7'd086, 7'd090}, '{7'd091, 7'd079, 7'd087, 7'd091}, '{7'd071, 7'd086, 7'd092, 7'd092}, '{7'd079, 7'd087, 7'd093, 7'd093}, '{7'd087, 7'd094, 7'd094, 7'd094}, '{7'd095, 7'd095, 7'd095, 7'd095},
      '{7'd096, 7'd096, 7'd096, 7'd096}, '{7'd104, 7'd097, 7'd097, 7'd097}, '{7'd112, 7'd104, 7'd098, 7'd098}, '{7'd120, 7'd105, 7'd099, 7'd099}, '{7'd100, 7'd112, 7'd104, 7'd100}, '{7'd108, 7'd113, 7'd105, 7'd101}, '{7'd116, 7'd120, 7'd106, 7'd102}, '{7'd124, 7'd121, 7'd107, 7'd103},
      '{7'd098, 7'd100, 7'd112, 7'd104}, '{7'd106, 7'd101, 7'd113, 7'd105}, '{7'd114, 7'd108, 7'd114, 7'd106}, '{7'd122, 7'd109, 7'd115, 7'd107}, '{7'd102, 7'd116, 7'd120, 7'd108}, '{7'd110, 7'd117, 7'd121, 7'd109}, '{7'd118, 7'd124, 7'd122, 7'd110}, '{7'd126, 7'd125, 7'd123, 7'd111},
      '{7'd097, 7'd098, 7'd100, 7'd112}, '{7'd105, 7'd099, 7'd101, 7'd113}, '{7'd113, 7'd106, 7'd102, 7'd114}, '{7'd121, 7'd107, 7'd103, 7'd115}, '{7'd101, 7'd114, 7'd108, 7'd116}, '{7'd109, 7'd115, 7'd109, 7'd117}, '{7'd117, 7'd122, 7'd110, 7'd118}, '{7'd125, 7'd123, 7'd111, 7'd119},
      '{7'd099, 7'd102, 7'd116, 7'd120}, '{7'd107, 7'd103, 7'd117, 7'd121}, '{7'd115, 7'd110, 7'd118, 7'd122}, '{7'd123, 7'd111, 7'd119, 7'd123}, '{7'd103, 7'd118, 7'd124, 7'd124}, '{7'd111, 7'd119, 7'd125, 7'd125}, '{7'd119, 7'd126, 7'd126, 7'd126}, '{7'd127, 7'd127, 7'd127, 7'd127}
    };

    automatic logic [8-1:0] lut_8lane [0:255][0:3] = '{
      '{8'd000, 8'd000, 8'd000, 8'd000}, '{8'd008, 8'd001, 8'd001, 8'd001}, '{8'd016, 8'd008, 8'd002, 8'd002}, '{8'd024, 8'd009, 8'd003, 8'd003}, '{8'd004, 8'd016, 8'd008, 8'd004}, '{8'd012, 8'd017, 8'd009, 8'd005}, '{8'd020, 8'd024, 8'd010, 8'd006}, '{8'd028, 8'd025, 8'd011, 8'd007},
      '{8'd002, 8'd004, 8'd016, 8'd008}, '{8'd010, 8'd005, 8'd017, 8'd009}, '{8'd018, 8'd012, 8'd018, 8'd010}, '{8'd026, 8'd013, 8'd019, 8'd011}, '{8'd006, 8'd020, 8'd024, 8'd012}, '{8'd014, 8'd021, 8'd025, 8'd013}, '{8'd022, 8'd028, 8'd026, 8'd014}, '{8'd030, 8'd029, 8'd027, 8'd015},
      '{8'd001, 8'd002, 8'd004, 8'd016}, '{8'd009, 8'd003, 8'd005, 8'd017}, '{8'd017, 8'd010, 8'd006, 8'd018}, '{8'd025, 8'd011, 8'd007, 8'd019}, '{8'd005, 8'd018, 8'd012, 8'd020}, '{8'd013, 8'd019, 8'd013, 8'd021}, '{8'd021, 8'd026, 8'd014, 8'd022}, '{8'd029, 8'd027, 8'd015, 8'd023},
      '{8'd003, 8'd006, 8'd020, 8'd024}, '{8'd011, 8'd007, 8'd021, 8'd025}, '{8'd019, 8'd014, 8'd022, 8'd026}, '{8'd027, 8'd015, 8'd023, 8'd027}, '{8'd007, 8'd022, 8'd028, 8'd028}, '{8'd015, 8'd023, 8'd029, 8'd029}, '{8'd023, 8'd030, 8'd030, 8'd030}, '{8'd031, 8'd031, 8'd031, 8'd031},
      '{8'd032, 8'd032, 8'd032, 8'd032}, '{8'd040, 8'd033, 8'd033, 8'd033}, '{8'd048, 8'd040, 8'd034, 8'd034}, '{8'd056, 8'd041, 8'd035, 8'd035}, '{8'd036, 8'd048, 8'd040, 8'd036}, '{8'd044, 8'd049, 8'd041, 8'd037}, '{8'd052, 8'd056, 8'd042, 8'd038}, '{8'd060, 8'd057, 8'd043, 8'd039},
      '{8'd034, 8'd036, 8'd048, 8'd040}, '{8'd042, 8'd037, 8'd049, 8'd041}, '{8'd050, 8'd044, 8'd050, 8'd042}, '{8'd058, 8'd045, 8'd051, 8'd043}, '{8'd038, 8'd052, 8'd056, 8'd044}, '{8'd046, 8'd053, 8'd057, 8'd045}, '{8'd054, 8'd060, 8'd058, 8'd046}, '{8'd062, 8'd061, 8'd059, 8'd047},
      '{8'd033, 8'd034, 8'd036, 8'd048}, '{8'd041, 8'd035, 8'd037, 8'd049}, '{8'd049, 8'd042, 8'd038, 8'd050}, '{8'd057, 8'd043, 8'd039, 8'd051}, '{8'd037, 8'd050, 8'd044, 8'd052}, '{8'd045, 8'd051, 8'd045, 8'd053}, '{8'd053, 8'd058, 8'd046, 8'd054}, '{8'd061, 8'd059, 8'd047, 8'd055},
      '{8'd035, 8'd038, 8'd052, 8'd056}, '{8'd043, 8'd039, 8'd053, 8'd057}, '{8'd051, 8'd046, 8'd054, 8'd058}, '{8'd059, 8'd047, 8'd055, 8'd059}, '{8'd039, 8'd054, 8'd060, 8'd060}, '{8'd047, 8'd055, 8'd061, 8'd061}, '{8'd055, 8'd062, 8'd062, 8'd062}, '{8'd063, 8'd063, 8'd063, 8'd063},
      '{8'd064, 8'd064, 8'd064, 8'd064}, '{8'd072, 8'd065, 8'd065, 8'd065}, '{8'd080, 8'd072, 8'd066, 8'd066}, '{8'd088, 8'd073, 8'd067, 8'd067}, '{8'd068, 8'd080, 8'd072, 8'd068}, '{8'd076, 8'd081, 8'd073, 8'd069}, '{8'd084, 8'd088, 8'd074, 8'd070}, '{8'd092, 8'd089, 8'd075, 8'd071},
      '{8'd066, 8'd068, 8'd080, 8'd072}, '{8'd074, 8'd069, 8'd081, 8'd073}, '{8'd082, 8'd076, 8'd082, 8'd074}, '{8'd090, 8'd077, 8'd083, 8'd075}, '{8'd070, 8'd084, 8'd088, 8'd076}, '{8'd078, 8'd085, 8'd089, 8'd077}, '{8'd086, 8'd092, 8'd090, 8'd078}, '{8'd094, 8'd093, 8'd091, 8'd079},
      '{8'd065, 8'd066, 8'd068, 8'd080}, '{8'd073, 8'd067, 8'd069, 8'd081}, '{8'd081, 8'd074, 8'd070, 8'd082}, '{8'd089, 8'd075, 8'd071, 8'd083}, '{8'd069, 8'd082, 8'd076, 8'd084}, '{8'd077, 8'd083, 8'd077, 8'd085}, '{8'd085, 8'd090, 8'd078, 8'd086}, '{8'd093, 8'd091, 8'd079, 8'd087},
      '{8'd067, 8'd070, 8'd084, 8'd088}, '{8'd075, 8'd071, 8'd085, 8'd089}, '{8'd083, 8'd078, 8'd086, 8'd090}, '{8'd091, 8'd079, 8'd087, 8'd091}, '{8'd071, 8'd086, 8'd092, 8'd092}, '{8'd079, 8'd087, 8'd093, 8'd093}, '{8'd087, 8'd094, 8'd094, 8'd094}, '{8'd095, 8'd095, 8'd095, 8'd095},
      '{8'd096, 8'd096, 8'd096, 8'd096}, '{8'd104, 8'd097, 8'd097, 8'd097}, '{8'd112, 8'd104, 8'd098, 8'd098}, '{8'd120, 8'd105, 8'd099, 8'd099}, '{8'd100, 8'd112, 8'd104, 8'd100}, '{8'd108, 8'd113, 8'd105, 8'd101}, '{8'd116, 8'd120, 8'd106, 8'd102}, '{8'd124, 8'd121, 8'd107, 8'd103},
      '{8'd098, 8'd100, 8'd112, 8'd104}, '{8'd106, 8'd101, 8'd113, 8'd105}, '{8'd114, 8'd108, 8'd114, 8'd106}, '{8'd122, 8'd109, 8'd115, 8'd107}, '{8'd102, 8'd116, 8'd120, 8'd108}, '{8'd110, 8'd117, 8'd121, 8'd109}, '{8'd118, 8'd124, 8'd122, 8'd110}, '{8'd126, 8'd125, 8'd123, 8'd111},
      '{8'd097, 8'd098, 8'd100, 8'd112}, '{8'd105, 8'd099, 8'd101, 8'd113}, '{8'd113, 8'd106, 8'd102, 8'd114}, '{8'd121, 8'd107, 8'd103, 8'd115}, '{8'd101, 8'd114, 8'd108, 8'd116}, '{8'd109, 8'd115, 8'd109, 8'd117}, '{8'd117, 8'd122, 8'd110, 8'd118}, '{8'd125, 8'd123, 8'd111, 8'd119},
      '{8'd099, 8'd102, 8'd116, 8'd120}, '{8'd107, 8'd103, 8'd117, 8'd121}, '{8'd115, 8'd110, 8'd118, 8'd122}, '{8'd123, 8'd111, 8'd119, 8'd123}, '{8'd103, 8'd118, 8'd124, 8'd124}, '{8'd111, 8'd119, 8'd125, 8'd125}, '{8'd119, 8'd126, 8'd126, 8'd126}, '{8'd127, 8'd127, 8'd127, 8'd127},
      '{8'd128, 8'd128, 8'd128, 8'd128}, '{8'd136, 8'd129, 8'd129, 8'd129}, '{8'd144, 8'd136, 8'd130, 8'd130}, '{8'd152, 8'd137, 8'd131, 8'd131}, '{8'd132, 8'd144, 8'd136, 8'd132}, '{8'd140, 8'd145, 8'd137, 8'd133}, '{8'd148, 8'd152, 8'd138, 8'd134}, '{8'd156, 8'd153, 8'd139, 8'd135},
      '{8'd130, 8'd132, 8'd144, 8'd136}, '{8'd138, 8'd133, 8'd145, 8'd137}, '{8'd146, 8'd140, 8'd146, 8'd138}, '{8'd154, 8'd141, 8'd147, 8'd139}, '{8'd134, 8'd148, 8'd152, 8'd140}, '{8'd142, 8'd149, 8'd153, 8'd141}, '{8'd150, 8'd156, 8'd154, 8'd142}, '{8'd158, 8'd157, 8'd155, 8'd143},
      '{8'd129, 8'd130, 8'd132, 8'd144}, '{8'd137, 8'd131, 8'd133, 8'd145}, '{8'd145, 8'd138, 8'd134, 8'd146}, '{8'd153, 8'd139, 8'd135, 8'd147}, '{8'd133, 8'd146, 8'd140, 8'd148}, '{8'd141, 8'd147, 8'd141, 8'd149}, '{8'd149, 8'd154, 8'd142, 8'd150}, '{8'd157, 8'd155, 8'd143, 8'd151},
      '{8'd131, 8'd134, 8'd148, 8'd152}, '{8'd139, 8'd135, 8'd149, 8'd153}, '{8'd147, 8'd142, 8'd150, 8'd154}, '{8'd155, 8'd143, 8'd151, 8'd155}, '{8'd135, 8'd150, 8'd156, 8'd156}, '{8'd143, 8'd151, 8'd157, 8'd157}, '{8'd151, 8'd158, 8'd158, 8'd158}, '{8'd159, 8'd159, 8'd159, 8'd159},
      '{8'd160, 8'd160, 8'd160, 8'd160}, '{8'd168, 8'd161, 8'd161, 8'd161}, '{8'd176, 8'd168, 8'd162, 8'd162}, '{8'd184, 8'd169, 8'd163, 8'd163}, '{8'd164, 8'd176, 8'd168, 8'd164}, '{8'd172, 8'd177, 8'd169, 8'd165}, '{8'd180, 8'd184, 8'd170, 8'd166}, '{8'd188, 8'd185, 8'd171, 8'd167},
      '{8'd162, 8'd164, 8'd176, 8'd168}, '{8'd170, 8'd165, 8'd177, 8'd169}, '{8'd178, 8'd172, 8'd178, 8'd170}, '{8'd186, 8'd173, 8'd179, 8'd171}, '{8'd166, 8'd180, 8'd184, 8'd172}, '{8'd174, 8'd181, 8'd185, 8'd173}, '{8'd182, 8'd188, 8'd186, 8'd174}, '{8'd190, 8'd189, 8'd187, 8'd175},
      '{8'd161, 8'd162, 8'd164, 8'd176}, '{8'd169, 8'd163, 8'd165, 8'd177}, '{8'd177, 8'd170, 8'd166, 8'd178}, '{8'd185, 8'd171, 8'd167, 8'd179}, '{8'd165, 8'd178, 8'd172, 8'd180}, '{8'd173, 8'd179, 8'd173, 8'd181}, '{8'd181, 8'd186, 8'd174, 8'd182}, '{8'd189, 8'd187, 8'd175, 8'd183},
      '{8'd163, 8'd166, 8'd180, 8'd184}, '{8'd171, 8'd167, 8'd181, 8'd185}, '{8'd179, 8'd174, 8'd182, 8'd186}, '{8'd187, 8'd175, 8'd183, 8'd187}, '{8'd167, 8'd182, 8'd188, 8'd188}, '{8'd175, 8'd183, 8'd189, 8'd189}, '{8'd183, 8'd190, 8'd190, 8'd190}, '{8'd191, 8'd191, 8'd191, 8'd191},
      '{8'd192, 8'd192, 8'd192, 8'd192}, '{8'd200, 8'd193, 8'd193, 8'd193}, '{8'd208, 8'd200, 8'd194, 8'd194}, '{8'd216, 8'd201, 8'd195, 8'd195}, '{8'd196, 8'd208, 8'd200, 8'd196}, '{8'd204, 8'd209, 8'd201, 8'd197}, '{8'd212, 8'd216, 8'd202, 8'd198}, '{8'd220, 8'd217, 8'd203, 8'd199},
      '{8'd194, 8'd196, 8'd208, 8'd200}, '{8'd202, 8'd197, 8'd209, 8'd201}, '{8'd210, 8'd204, 8'd210, 8'd202}, '{8'd218, 8'd205, 8'd211, 8'd203}, '{8'd198, 8'd212, 8'd216, 8'd204}, '{8'd206, 8'd213, 8'd217, 8'd205}, '{8'd214, 8'd220, 8'd218, 8'd206}, '{8'd222, 8'd221, 8'd219, 8'd207},
      '{8'd193, 8'd194, 8'd196, 8'd208}, '{8'd201, 8'd195, 8'd197, 8'd209}, '{8'd209, 8'd202, 8'd198, 8'd210}, '{8'd217, 8'd203, 8'd199, 8'd211}, '{8'd197, 8'd210, 8'd204, 8'd212}, '{8'd205, 8'd211, 8'd205, 8'd213}, '{8'd213, 8'd218, 8'd206, 8'd214}, '{8'd221, 8'd219, 8'd207, 8'd215},
      '{8'd195, 8'd198, 8'd212, 8'd216}, '{8'd203, 8'd199, 8'd213, 8'd217}, '{8'd211, 8'd206, 8'd214, 8'd218}, '{8'd219, 8'd207, 8'd215, 8'd219}, '{8'd199, 8'd214, 8'd220, 8'd220}, '{8'd207, 8'd215, 8'd221, 8'd221}, '{8'd215, 8'd222, 8'd222, 8'd222}, '{8'd223, 8'd223, 8'd223, 8'd223},
      '{8'd224, 8'd224, 8'd224, 8'd224}, '{8'd232, 8'd225, 8'd225, 8'd225}, '{8'd240, 8'd232, 8'd226, 8'd226}, '{8'd248, 8'd233, 8'd227, 8'd227}, '{8'd228, 8'd240, 8'd232, 8'd228}, '{8'd236, 8'd241, 8'd233, 8'd229}, '{8'd244, 8'd248, 8'd234, 8'd230}, '{8'd252, 8'd249, 8'd235, 8'd231},
      '{8'd226, 8'd228, 8'd240, 8'd232}, '{8'd234, 8'd229, 8'd241, 8'd233}, '{8'd242, 8'd236, 8'd242, 8'd234}, '{8'd250, 8'd237, 8'd243, 8'd235}, '{8'd230, 8'd244, 8'd248, 8'd236}, '{8'd238, 8'd245, 8'd249, 8'd237}, '{8'd246, 8'd252, 8'd250, 8'd238}, '{8'd254, 8'd253, 8'd251, 8'd239},
      '{8'd225, 8'd226, 8'd228, 8'd240}, '{8'd233, 8'd227, 8'd229, 8'd241}, '{8'd241, 8'd234, 8'd230, 8'd242}, '{8'd249, 8'd235, 8'd231, 8'd243}, '{8'd229, 8'd242, 8'd236, 8'd244}, '{8'd237, 8'd243, 8'd237, 8'd245}, '{8'd245, 8'd250, 8'd238, 8'd246}, '{8'd253, 8'd251, 8'd239, 8'd247},
      '{8'd227, 8'd230, 8'd244, 8'd248}, '{8'd235, 8'd231, 8'd245, 8'd249}, '{8'd243, 8'd238, 8'd246, 8'd250}, '{8'd251, 8'd239, 8'd247, 8'd251}, '{8'd231, 8'd246, 8'd252, 8'd252}, '{8'd239, 8'd247, 8'd253, 8'd253}, '{8'd247, 8'd254, 8'd254, 8'd254}, '{8'd255, 8'd255, 8'd255, 8'd255}
    };

    automatic logic [9-1:0] lut_16lane [0:511][0:3] = '{
      '{9'd000, 9'd000, 9'd000, 9'd000}, '{9'd008, 9'd001, 9'd001, 9'd001}, '{9'd016, 9'd008, 9'd002, 9'd002}, '{9'd024, 9'd009, 9'd003, 9'd003}, '{9'd004, 9'd016, 9'd008, 9'd004}, '{9'd012, 9'd017, 9'd009, 9'd005}, '{9'd020, 9'd024, 9'd010, 9'd006}, '{9'd028, 9'd025, 9'd011, 9'd007},
      '{9'd002, 9'd004, 9'd016, 9'd008}, '{9'd010, 9'd005, 9'd017, 9'd009}, '{9'd018, 9'd012, 9'd018, 9'd010}, '{9'd026, 9'd013, 9'd019, 9'd011}, '{9'd006, 9'd020, 9'd024, 9'd012}, '{9'd014, 9'd021, 9'd025, 9'd013}, '{9'd022, 9'd028, 9'd026, 9'd014}, '{9'd030, 9'd029, 9'd027, 9'd015},
      '{9'd001, 9'd002, 9'd004, 9'd016}, '{9'd009, 9'd003, 9'd005, 9'd017}, '{9'd017, 9'd010, 9'd006, 9'd018}, '{9'd025, 9'd011, 9'd007, 9'd019}, '{9'd005, 9'd018, 9'd012, 9'd020}, '{9'd013, 9'd019, 9'd013, 9'd021}, '{9'd021, 9'd026, 9'd014, 9'd022}, '{9'd029, 9'd027, 9'd015, 9'd023},
      '{9'd003, 9'd006, 9'd020, 9'd024}, '{9'd011, 9'd007, 9'd021, 9'd025}, '{9'd019, 9'd014, 9'd022, 9'd026}, '{9'd027, 9'd015, 9'd023, 9'd027}, '{9'd007, 9'd022, 9'd028, 9'd028}, '{9'd015, 9'd023, 9'd029, 9'd029}, '{9'd023, 9'd030, 9'd030, 9'd030}, '{9'd031, 9'd031, 9'd031, 9'd031},
      '{9'd032, 9'd032, 9'd032, 9'd032}, '{9'd040, 9'd033, 9'd033, 9'd033}, '{9'd048, 9'd040, 9'd034, 9'd034}, '{9'd056, 9'd041, 9'd035, 9'd035}, '{9'd036, 9'd048, 9'd040, 9'd036}, '{9'd044, 9'd049, 9'd041, 9'd037}, '{9'd052, 9'd056, 9'd042, 9'd038}, '{9'd060, 9'd057, 9'd043, 9'd039},
      '{9'd034, 9'd036, 9'd048, 9'd040}, '{9'd042, 9'd037, 9'd049, 9'd041}, '{9'd050, 9'd044, 9'd050, 9'd042}, '{9'd058, 9'd045, 9'd051, 9'd043}, '{9'd038, 9'd052, 9'd056, 9'd044}, '{9'd046, 9'd053, 9'd057, 9'd045}, '{9'd054, 9'd060, 9'd058, 9'd046}, '{9'd062, 9'd061, 9'd059, 9'd047},
      '{9'd033, 9'd034, 9'd036, 9'd048}, '{9'd041, 9'd035, 9'd037, 9'd049}, '{9'd049, 9'd042, 9'd038, 9'd050}, '{9'd057, 9'd043, 9'd039, 9'd051}, '{9'd037, 9'd050, 9'd044, 9'd052}, '{9'd045, 9'd051, 9'd045, 9'd053}, '{9'd053, 9'd058, 9'd046, 9'd054}, '{9'd061, 9'd059, 9'd047, 9'd055},
      '{9'd035, 9'd038, 9'd052, 9'd056}, '{9'd043, 9'd039, 9'd053, 9'd057}, '{9'd051, 9'd046, 9'd054, 9'd058}, '{9'd059, 9'd047, 9'd055, 9'd059}, '{9'd039, 9'd054, 9'd060, 9'd060}, '{9'd047, 9'd055, 9'd061, 9'd061}, '{9'd055, 9'd062, 9'd062, 9'd062}, '{9'd063, 9'd063, 9'd063, 9'd063},
      '{9'd064, 9'd064, 9'd064, 9'd064}, '{9'd072, 9'd065, 9'd065, 9'd065}, '{9'd080, 9'd072, 9'd066, 9'd066}, '{9'd088, 9'd073, 9'd067, 9'd067}, '{9'd068, 9'd080, 9'd072, 9'd068}, '{9'd076, 9'd081, 9'd073, 9'd069}, '{9'd084, 9'd088, 9'd074, 9'd070}, '{9'd092, 9'd089, 9'd075, 9'd071},
      '{9'd066, 9'd068, 9'd080, 9'd072}, '{9'd074, 9'd069, 9'd081, 9'd073}, '{9'd082, 9'd076, 9'd082, 9'd074}, '{9'd090, 9'd077, 9'd083, 9'd075}, '{9'd070, 9'd084, 9'd088, 9'd076}, '{9'd078, 9'd085, 9'd089, 9'd077}, '{9'd086, 9'd092, 9'd090, 9'd078}, '{9'd094, 9'd093, 9'd091, 9'd079},
      '{9'd065, 9'd066, 9'd068, 9'd080}, '{9'd073, 9'd067, 9'd069, 9'd081}, '{9'd081, 9'd074, 9'd070, 9'd082}, '{9'd089, 9'd075, 9'd071, 9'd083}, '{9'd069, 9'd082, 9'd076, 9'd084}, '{9'd077, 9'd083, 9'd077, 9'd085}, '{9'd085, 9'd090, 9'd078, 9'd086}, '{9'd093, 9'd091, 9'd079, 9'd087},
      '{9'd067, 9'd070, 9'd084, 9'd088}, '{9'd075, 9'd071, 9'd085, 9'd089}, '{9'd083, 9'd078, 9'd086, 9'd090}, '{9'd091, 9'd079, 9'd087, 9'd091}, '{9'd071, 9'd086, 9'd092, 9'd092}, '{9'd079, 9'd087, 9'd093, 9'd093}, '{9'd087, 9'd094, 9'd094, 9'd094}, '{9'd095, 9'd095, 9'd095, 9'd095},
      '{9'd096, 9'd096, 9'd096, 9'd096}, '{9'd104, 9'd097, 9'd097, 9'd097}, '{9'd112, 9'd104, 9'd098, 9'd098}, '{9'd120, 9'd105, 9'd099, 9'd099}, '{9'd100, 9'd112, 9'd104, 9'd100}, '{9'd108, 9'd113, 9'd105, 9'd101}, '{9'd116, 9'd120, 9'd106, 9'd102}, '{9'd124, 9'd121, 9'd107, 9'd103},
      '{9'd098, 9'd100, 9'd112, 9'd104}, '{9'd106, 9'd101, 9'd113, 9'd105}, '{9'd114, 9'd108, 9'd114, 9'd106}, '{9'd122, 9'd109, 9'd115, 9'd107}, '{9'd102, 9'd116, 9'd120, 9'd108}, '{9'd110, 9'd117, 9'd121, 9'd109}, '{9'd118, 9'd124, 9'd122, 9'd110}, '{9'd126, 9'd125, 9'd123, 9'd111},
      '{9'd097, 9'd098, 9'd100, 9'd112}, '{9'd105, 9'd099, 9'd101, 9'd113}, '{9'd113, 9'd106, 9'd102, 9'd114}, '{9'd121, 9'd107, 9'd103, 9'd115}, '{9'd101, 9'd114, 9'd108, 9'd116}, '{9'd109, 9'd115, 9'd109, 9'd117}, '{9'd117, 9'd122, 9'd110, 9'd118}, '{9'd125, 9'd123, 9'd111, 9'd119},
      '{9'd099, 9'd102, 9'd116, 9'd120}, '{9'd107, 9'd103, 9'd117, 9'd121}, '{9'd115, 9'd110, 9'd118, 9'd122}, '{9'd123, 9'd111, 9'd119, 9'd123}, '{9'd103, 9'd118, 9'd124, 9'd124}, '{9'd111, 9'd119, 9'd125, 9'd125}, '{9'd119, 9'd126, 9'd126, 9'd126}, '{9'd127, 9'd127, 9'd127, 9'd127},
      '{9'd128, 9'd128, 9'd128, 9'd128}, '{9'd136, 9'd129, 9'd129, 9'd129}, '{9'd144, 9'd136, 9'd130, 9'd130}, '{9'd152, 9'd137, 9'd131, 9'd131}, '{9'd132, 9'd144, 9'd136, 9'd132}, '{9'd140, 9'd145, 9'd137, 9'd133}, '{9'd148, 9'd152, 9'd138, 9'd134}, '{9'd156, 9'd153, 9'd139, 9'd135},
      '{9'd130, 9'd132, 9'd144, 9'd136}, '{9'd138, 9'd133, 9'd145, 9'd137}, '{9'd146, 9'd140, 9'd146, 9'd138}, '{9'd154, 9'd141, 9'd147, 9'd139}, '{9'd134, 9'd148, 9'd152, 9'd140}, '{9'd142, 9'd149, 9'd153, 9'd141}, '{9'd150, 9'd156, 9'd154, 9'd142}, '{9'd158, 9'd157, 9'd155, 9'd143},
      '{9'd129, 9'd130, 9'd132, 9'd144}, '{9'd137, 9'd131, 9'd133, 9'd145}, '{9'd145, 9'd138, 9'd134, 9'd146}, '{9'd153, 9'd139, 9'd135, 9'd147}, '{9'd133, 9'd146, 9'd140, 9'd148}, '{9'd141, 9'd147, 9'd141, 9'd149}, '{9'd149, 9'd154, 9'd142, 9'd150}, '{9'd157, 9'd155, 9'd143, 9'd151},
      '{9'd131, 9'd134, 9'd148, 9'd152}, '{9'd139, 9'd135, 9'd149, 9'd153}, '{9'd147, 9'd142, 9'd150, 9'd154}, '{9'd155, 9'd143, 9'd151, 9'd155}, '{9'd135, 9'd150, 9'd156, 9'd156}, '{9'd143, 9'd151, 9'd157, 9'd157}, '{9'd151, 9'd158, 9'd158, 9'd158}, '{9'd159, 9'd159, 9'd159, 9'd159},
      '{9'd160, 9'd160, 9'd160, 9'd160}, '{9'd168, 9'd161, 9'd161, 9'd161}, '{9'd176, 9'd168, 9'd162, 9'd162}, '{9'd184, 9'd169, 9'd163, 9'd163}, '{9'd164, 9'd176, 9'd168, 9'd164}, '{9'd172, 9'd177, 9'd169, 9'd165}, '{9'd180, 9'd184, 9'd170, 9'd166}, '{9'd188, 9'd185, 9'd171, 9'd167},
      '{9'd162, 9'd164, 9'd176, 9'd168}, '{9'd170, 9'd165, 9'd177, 9'd169}, '{9'd178, 9'd172, 9'd178, 9'd170}, '{9'd186, 9'd173, 9'd179, 9'd171}, '{9'd166, 9'd180, 9'd184, 9'd172}, '{9'd174, 9'd181, 9'd185, 9'd173}, '{9'd182, 9'd188, 9'd186, 9'd174}, '{9'd190, 9'd189, 9'd187, 9'd175},
      '{9'd161, 9'd162, 9'd164, 9'd176}, '{9'd169, 9'd163, 9'd165, 9'd177}, '{9'd177, 9'd170, 9'd166, 9'd178}, '{9'd185, 9'd171, 9'd167, 9'd179}, '{9'd165, 9'd178, 9'd172, 9'd180}, '{9'd173, 9'd179, 9'd173, 9'd181}, '{9'd181, 9'd186, 9'd174, 9'd182}, '{9'd189, 9'd187, 9'd175, 9'd183},
      '{9'd163, 9'd166, 9'd180, 9'd184}, '{9'd171, 9'd167, 9'd181, 9'd185}, '{9'd179, 9'd174, 9'd182, 9'd186}, '{9'd187, 9'd175, 9'd183, 9'd187}, '{9'd167, 9'd182, 9'd188, 9'd188}, '{9'd175, 9'd183, 9'd189, 9'd189}, '{9'd183, 9'd190, 9'd190, 9'd190}, '{9'd191, 9'd191, 9'd191, 9'd191},
      '{9'd192, 9'd192, 9'd192, 9'd192}, '{9'd200, 9'd193, 9'd193, 9'd193}, '{9'd208, 9'd200, 9'd194, 9'd194}, '{9'd216, 9'd201, 9'd195, 9'd195}, '{9'd196, 9'd208, 9'd200, 9'd196}, '{9'd204, 9'd209, 9'd201, 9'd197}, '{9'd212, 9'd216, 9'd202, 9'd198}, '{9'd220, 9'd217, 9'd203, 9'd199},
      '{9'd194, 9'd196, 9'd208, 9'd200}, '{9'd202, 9'd197, 9'd209, 9'd201}, '{9'd210, 9'd204, 9'd210, 9'd202}, '{9'd218, 9'd205, 9'd211, 9'd203}, '{9'd198, 9'd212, 9'd216, 9'd204}, '{9'd206, 9'd213, 9'd217, 9'd205}, '{9'd214, 9'd220, 9'd218, 9'd206}, '{9'd222, 9'd221, 9'd219, 9'd207},
      '{9'd193, 9'd194, 9'd196, 9'd208}, '{9'd201, 9'd195, 9'd197, 9'd209}, '{9'd209, 9'd202, 9'd198, 9'd210}, '{9'd217, 9'd203, 9'd199, 9'd211}, '{9'd197, 9'd210, 9'd204, 9'd212}, '{9'd205, 9'd211, 9'd205, 9'd213}, '{9'd213, 9'd218, 9'd206, 9'd214}, '{9'd221, 9'd219, 9'd207, 9'd215},
      '{9'd195, 9'd198, 9'd212, 9'd216}, '{9'd203, 9'd199, 9'd213, 9'd217}, '{9'd211, 9'd206, 9'd214, 9'd218}, '{9'd219, 9'd207, 9'd215, 9'd219}, '{9'd199, 9'd214, 9'd220, 9'd220}, '{9'd207, 9'd215, 9'd221, 9'd221}, '{9'd215, 9'd222, 9'd222, 9'd222}, '{9'd223, 9'd223, 9'd223, 9'd223},
      '{9'd224, 9'd224, 9'd224, 9'd224}, '{9'd232, 9'd225, 9'd225, 9'd225}, '{9'd240, 9'd232, 9'd226, 9'd226}, '{9'd248, 9'd233, 9'd227, 9'd227}, '{9'd228, 9'd240, 9'd232, 9'd228}, '{9'd236, 9'd241, 9'd233, 9'd229}, '{9'd244, 9'd248, 9'd234, 9'd230}, '{9'd252, 9'd249, 9'd235, 9'd231},
      '{9'd226, 9'd228, 9'd240, 9'd232}, '{9'd234, 9'd229, 9'd241, 9'd233}, '{9'd242, 9'd236, 9'd242, 9'd234}, '{9'd250, 9'd237, 9'd243, 9'd235}, '{9'd230, 9'd244, 9'd248, 9'd236}, '{9'd238, 9'd245, 9'd249, 9'd237}, '{9'd246, 9'd252, 9'd250, 9'd238}, '{9'd254, 9'd253, 9'd251, 9'd239},
      '{9'd225, 9'd226, 9'd228, 9'd240}, '{9'd233, 9'd227, 9'd229, 9'd241}, '{9'd241, 9'd234, 9'd230, 9'd242}, '{9'd249, 9'd235, 9'd231, 9'd243}, '{9'd229, 9'd242, 9'd236, 9'd244}, '{9'd237, 9'd243, 9'd237, 9'd245}, '{9'd245, 9'd250, 9'd238, 9'd246}, '{9'd253, 9'd251, 9'd239, 9'd247},
      '{9'd227, 9'd230, 9'd244, 9'd248}, '{9'd235, 9'd231, 9'd245, 9'd249}, '{9'd243, 9'd238, 9'd246, 9'd250}, '{9'd251, 9'd239, 9'd247, 9'd251}, '{9'd231, 9'd246, 9'd252, 9'd252}, '{9'd239, 9'd247, 9'd253, 9'd253}, '{9'd247, 9'd254, 9'd254, 9'd254}, '{9'd255, 9'd255, 9'd255, 9'd255},
      '{9'd256, 9'd256, 9'd256, 9'd256}, '{9'd264, 9'd257, 9'd257, 9'd257}, '{9'd272, 9'd264, 9'd258, 9'd258}, '{9'd280, 9'd265, 9'd259, 9'd259}, '{9'd260, 9'd272, 9'd264, 9'd260}, '{9'd268, 9'd273, 9'd265, 9'd261}, '{9'd276, 9'd280, 9'd266, 9'd262}, '{9'd284, 9'd281, 9'd267, 9'd263},
      '{9'd258, 9'd260, 9'd272, 9'd264}, '{9'd266, 9'd261, 9'd273, 9'd265}, '{9'd274, 9'd268, 9'd274, 9'd266}, '{9'd282, 9'd269, 9'd275, 9'd267}, '{9'd262, 9'd276, 9'd280, 9'd268}, '{9'd270, 9'd277, 9'd281, 9'd269}, '{9'd278, 9'd284, 9'd282, 9'd270}, '{9'd286, 9'd285, 9'd283, 9'd271},
      '{9'd257, 9'd258, 9'd260, 9'd272}, '{9'd265, 9'd259, 9'd261, 9'd273}, '{9'd273, 9'd266, 9'd262, 9'd274}, '{9'd281, 9'd267, 9'd263, 9'd275}, '{9'd261, 9'd274, 9'd268, 9'd276}, '{9'd269, 9'd275, 9'd269, 9'd277}, '{9'd277, 9'd282, 9'd270, 9'd278}, '{9'd285, 9'd283, 9'd271, 9'd279},
      '{9'd259, 9'd262, 9'd276, 9'd280}, '{9'd267, 9'd263, 9'd277, 9'd281}, '{9'd275, 9'd270, 9'd278, 9'd282}, '{9'd283, 9'd271, 9'd279, 9'd283}, '{9'd263, 9'd278, 9'd284, 9'd284}, '{9'd271, 9'd279, 9'd285, 9'd285}, '{9'd279, 9'd286, 9'd286, 9'd286}, '{9'd287, 9'd287, 9'd287, 9'd287},
      '{9'd288, 9'd288, 9'd288, 9'd288}, '{9'd296, 9'd289, 9'd289, 9'd289}, '{9'd304, 9'd296, 9'd290, 9'd290}, '{9'd312, 9'd297, 9'd291, 9'd291}, '{9'd292, 9'd304, 9'd296, 9'd292}, '{9'd300, 9'd305, 9'd297, 9'd293}, '{9'd308, 9'd312, 9'd298, 9'd294}, '{9'd316, 9'd313, 9'd299, 9'd295},
      '{9'd290, 9'd292, 9'd304, 9'd296}, '{9'd298, 9'd293, 9'd305, 9'd297}, '{9'd306, 9'd300, 9'd306, 9'd298}, '{9'd314, 9'd301, 9'd307, 9'd299}, '{9'd294, 9'd308, 9'd312, 9'd300}, '{9'd302, 9'd309, 9'd313, 9'd301}, '{9'd310, 9'd316, 9'd314, 9'd302}, '{9'd318, 9'd317, 9'd315, 9'd303},
      '{9'd289, 9'd290, 9'd292, 9'd304}, '{9'd297, 9'd291, 9'd293, 9'd305}, '{9'd305, 9'd298, 9'd294, 9'd306}, '{9'd313, 9'd299, 9'd295, 9'd307}, '{9'd293, 9'd306, 9'd300, 9'd308}, '{9'd301, 9'd307, 9'd301, 9'd309}, '{9'd309, 9'd314, 9'd302, 9'd310}, '{9'd317, 9'd315, 9'd303, 9'd311},
      '{9'd291, 9'd294, 9'd308, 9'd312}, '{9'd299, 9'd295, 9'd309, 9'd313}, '{9'd307, 9'd302, 9'd310, 9'd314}, '{9'd315, 9'd303, 9'd311, 9'd315}, '{9'd295, 9'd310, 9'd316, 9'd316}, '{9'd303, 9'd311, 9'd317, 9'd317}, '{9'd311, 9'd318, 9'd318, 9'd318}, '{9'd319, 9'd319, 9'd319, 9'd319},
      '{9'd320, 9'd320, 9'd320, 9'd320}, '{9'd328, 9'd321, 9'd321, 9'd321}, '{9'd336, 9'd328, 9'd322, 9'd322}, '{9'd344, 9'd329, 9'd323, 9'd323}, '{9'd324, 9'd336, 9'd328, 9'd324}, '{9'd332, 9'd337, 9'd329, 9'd325}, '{9'd340, 9'd344, 9'd330, 9'd326}, '{9'd348, 9'd345, 9'd331, 9'd327},
      '{9'd322, 9'd324, 9'd336, 9'd328}, '{9'd330, 9'd325, 9'd337, 9'd329}, '{9'd338, 9'd332, 9'd338, 9'd330}, '{9'd346, 9'd333, 9'd339, 9'd331}, '{9'd326, 9'd340, 9'd344, 9'd332}, '{9'd334, 9'd341, 9'd345, 9'd333}, '{9'd342, 9'd348, 9'd346, 9'd334}, '{9'd350, 9'd349, 9'd347, 9'd335},
      '{9'd321, 9'd322, 9'd324, 9'd336}, '{9'd329, 9'd323, 9'd325, 9'd337}, '{9'd337, 9'd330, 9'd326, 9'd338}, '{9'd345, 9'd331, 9'd327, 9'd339}, '{9'd325, 9'd338, 9'd332, 9'd340}, '{9'd333, 9'd339, 9'd333, 9'd341}, '{9'd341, 9'd346, 9'd334, 9'd342}, '{9'd349, 9'd347, 9'd335, 9'd343},
      '{9'd323, 9'd326, 9'd340, 9'd344}, '{9'd331, 9'd327, 9'd341, 9'd345}, '{9'd339, 9'd334, 9'd342, 9'd346}, '{9'd347, 9'd335, 9'd343, 9'd347}, '{9'd327, 9'd342, 9'd348, 9'd348}, '{9'd335, 9'd343, 9'd349, 9'd349}, '{9'd343, 9'd350, 9'd350, 9'd350}, '{9'd351, 9'd351, 9'd351, 9'd351},
      '{9'd352, 9'd352, 9'd352, 9'd352}, '{9'd360, 9'd353, 9'd353, 9'd353}, '{9'd368, 9'd360, 9'd354, 9'd354}, '{9'd376, 9'd361, 9'd355, 9'd355}, '{9'd356, 9'd368, 9'd360, 9'd356}, '{9'd364, 9'd369, 9'd361, 9'd357}, '{9'd372, 9'd376, 9'd362, 9'd358}, '{9'd380, 9'd377, 9'd363, 9'd359},
      '{9'd354, 9'd356, 9'd368, 9'd360}, '{9'd362, 9'd357, 9'd369, 9'd361}, '{9'd370, 9'd364, 9'd370, 9'd362}, '{9'd378, 9'd365, 9'd371, 9'd363}, '{9'd358, 9'd372, 9'd376, 9'd364}, '{9'd366, 9'd373, 9'd377, 9'd365}, '{9'd374, 9'd380, 9'd378, 9'd366}, '{9'd382, 9'd381, 9'd379, 9'd367},
      '{9'd353, 9'd354, 9'd356, 9'd368}, '{9'd361, 9'd355, 9'd357, 9'd369}, '{9'd369, 9'd362, 9'd358, 9'd370}, '{9'd377, 9'd363, 9'd359, 9'd371}, '{9'd357, 9'd370, 9'd364, 9'd372}, '{9'd365, 9'd371, 9'd365, 9'd373}, '{9'd373, 9'd378, 9'd366, 9'd374}, '{9'd381, 9'd379, 9'd367, 9'd375},
      '{9'd355, 9'd358, 9'd372, 9'd376}, '{9'd363, 9'd359, 9'd373, 9'd377}, '{9'd371, 9'd366, 9'd374, 9'd378}, '{9'd379, 9'd367, 9'd375, 9'd379}, '{9'd359, 9'd374, 9'd380, 9'd380}, '{9'd367, 9'd375, 9'd381, 9'd381}, '{9'd375, 9'd382, 9'd382, 9'd382}, '{9'd383, 9'd383, 9'd383, 9'd383},
      '{9'd384, 9'd384, 9'd384, 9'd384}, '{9'd392, 9'd385, 9'd385, 9'd385}, '{9'd400, 9'd392, 9'd386, 9'd386}, '{9'd408, 9'd393, 9'd387, 9'd387}, '{9'd388, 9'd400, 9'd392, 9'd388}, '{9'd396, 9'd401, 9'd393, 9'd389}, '{9'd404, 9'd408, 9'd394, 9'd390}, '{9'd412, 9'd409, 9'd395, 9'd391},
      '{9'd386, 9'd388, 9'd400, 9'd392}, '{9'd394, 9'd389, 9'd401, 9'd393}, '{9'd402, 9'd396, 9'd402, 9'd394}, '{9'd410, 9'd397, 9'd403, 9'd395}, '{9'd390, 9'd404, 9'd408, 9'd396}, '{9'd398, 9'd405, 9'd409, 9'd397}, '{9'd406, 9'd412, 9'd410, 9'd398}, '{9'd414, 9'd413, 9'd411, 9'd399},
      '{9'd385, 9'd386, 9'd388, 9'd400}, '{9'd393, 9'd387, 9'd389, 9'd401}, '{9'd401, 9'd394, 9'd390, 9'd402}, '{9'd409, 9'd395, 9'd391, 9'd403}, '{9'd389, 9'd402, 9'd396, 9'd404}, '{9'd397, 9'd403, 9'd397, 9'd405}, '{9'd405, 9'd410, 9'd398, 9'd406}, '{9'd413, 9'd411, 9'd399, 9'd407},
      '{9'd387, 9'd390, 9'd404, 9'd408}, '{9'd395, 9'd391, 9'd405, 9'd409}, '{9'd403, 9'd398, 9'd406, 9'd410}, '{9'd411, 9'd399, 9'd407, 9'd411}, '{9'd391, 9'd406, 9'd412, 9'd412}, '{9'd399, 9'd407, 9'd413, 9'd413}, '{9'd407, 9'd414, 9'd414, 9'd414}, '{9'd415, 9'd415, 9'd415, 9'd415},
      '{9'd416, 9'd416, 9'd416, 9'd416}, '{9'd424, 9'd417, 9'd417, 9'd417}, '{9'd432, 9'd424, 9'd418, 9'd418}, '{9'd440, 9'd425, 9'd419, 9'd419}, '{9'd420, 9'd432, 9'd424, 9'd420}, '{9'd428, 9'd433, 9'd425, 9'd421}, '{9'd436, 9'd440, 9'd426, 9'd422}, '{9'd444, 9'd441, 9'd427, 9'd423},
      '{9'd418, 9'd420, 9'd432, 9'd424}, '{9'd426, 9'd421, 9'd433, 9'd425}, '{9'd434, 9'd428, 9'd434, 9'd426}, '{9'd442, 9'd429, 9'd435, 9'd427}, '{9'd422, 9'd436, 9'd440, 9'd428}, '{9'd430, 9'd437, 9'd441, 9'd429}, '{9'd438, 9'd444, 9'd442, 9'd430}, '{9'd446, 9'd445, 9'd443, 9'd431},
      '{9'd417, 9'd418, 9'd420, 9'd432}, '{9'd425, 9'd419, 9'd421, 9'd433}, '{9'd433, 9'd426, 9'd422, 9'd434}, '{9'd441, 9'd427, 9'd423, 9'd435}, '{9'd421, 9'd434, 9'd428, 9'd436}, '{9'd429, 9'd435, 9'd429, 9'd437}, '{9'd437, 9'd442, 9'd430, 9'd438}, '{9'd445, 9'd443, 9'd431, 9'd439},
      '{9'd419, 9'd422, 9'd436, 9'd440}, '{9'd427, 9'd423, 9'd437, 9'd441}, '{9'd435, 9'd430, 9'd438, 9'd442}, '{9'd443, 9'd431, 9'd439, 9'd443}, '{9'd423, 9'd438, 9'd444, 9'd444}, '{9'd431, 9'd439, 9'd445, 9'd445}, '{9'd439, 9'd446, 9'd446, 9'd446}, '{9'd447, 9'd447, 9'd447, 9'd447},
      '{9'd448, 9'd448, 9'd448, 9'd448}, '{9'd456, 9'd449, 9'd449, 9'd449}, '{9'd464, 9'd456, 9'd450, 9'd450}, '{9'd472, 9'd457, 9'd451, 9'd451}, '{9'd452, 9'd464, 9'd456, 9'd452}, '{9'd460, 9'd465, 9'd457, 9'd453}, '{9'd468, 9'd472, 9'd458, 9'd454}, '{9'd476, 9'd473, 9'd459, 9'd455},
      '{9'd450, 9'd452, 9'd464, 9'd456}, '{9'd458, 9'd453, 9'd465, 9'd457}, '{9'd466, 9'd460, 9'd466, 9'd458}, '{9'd474, 9'd461, 9'd467, 9'd459}, '{9'd454, 9'd468, 9'd472, 9'd460}, '{9'd462, 9'd469, 9'd473, 9'd461}, '{9'd470, 9'd476, 9'd474, 9'd462}, '{9'd478, 9'd477, 9'd475, 9'd463},
      '{9'd449, 9'd450, 9'd452, 9'd464}, '{9'd457, 9'd451, 9'd453, 9'd465}, '{9'd465, 9'd458, 9'd454, 9'd466}, '{9'd473, 9'd459, 9'd455, 9'd467}, '{9'd453, 9'd466, 9'd460, 9'd468}, '{9'd461, 9'd467, 9'd461, 9'd469}, '{9'd469, 9'd474, 9'd462, 9'd470}, '{9'd477, 9'd475, 9'd463, 9'd471},
      '{9'd451, 9'd454, 9'd468, 9'd472}, '{9'd459, 9'd455, 9'd469, 9'd473}, '{9'd467, 9'd462, 9'd470, 9'd474}, '{9'd475, 9'd463, 9'd471, 9'd475}, '{9'd455, 9'd470, 9'd476, 9'd476}, '{9'd463, 9'd471, 9'd477, 9'd477}, '{9'd471, 9'd478, 9'd478, 9'd478}, '{9'd479, 9'd479, 9'd479, 9'd479},
      '{9'd480, 9'd480, 9'd480, 9'd480}, '{9'd488, 9'd481, 9'd481, 9'd481}, '{9'd496, 9'd488, 9'd482, 9'd482}, '{9'd504, 9'd489, 9'd483, 9'd483}, '{9'd484, 9'd496, 9'd488, 9'd484}, '{9'd492, 9'd497, 9'd489, 9'd485}, '{9'd500, 9'd504, 9'd490, 9'd486}, '{9'd508, 9'd505, 9'd491, 9'd487},
      '{9'd482, 9'd484, 9'd496, 9'd488}, '{9'd490, 9'd485, 9'd497, 9'd489}, '{9'd498, 9'd492, 9'd498, 9'd490}, '{9'd506, 9'd493, 9'd499, 9'd491}, '{9'd486, 9'd500, 9'd504, 9'd492}, '{9'd494, 9'd501, 9'd505, 9'd493}, '{9'd502, 9'd508, 9'd506, 9'd494}, '{9'd510, 9'd509, 9'd507, 9'd495},
      '{9'd481, 9'd482, 9'd484, 9'd496}, '{9'd489, 9'd483, 9'd485, 9'd497}, '{9'd497, 9'd490, 9'd486, 9'd498}, '{9'd505, 9'd491, 9'd487, 9'd499}, '{9'd485, 9'd498, 9'd492, 9'd500}, '{9'd493, 9'd499, 9'd493, 9'd501}, '{9'd501, 9'd506, 9'd494, 9'd502}, '{9'd509, 9'd507, 9'd495, 9'd503},
      '{9'd483, 9'd486, 9'd500, 9'd504}, '{9'd491, 9'd487, 9'd501, 9'd505}, '{9'd499, 9'd494, 9'd502, 9'd506}, '{9'd507, 9'd495, 9'd503, 9'd507}, '{9'd487, 9'd502, 9'd508, 9'd508}, '{9'd495, 9'd503, 9'd509, 9'd509}, '{9'd503, 9'd510, 9'd510, 9'd510}, '{9'd511, 9'd511, 9'd511, 9'd511}
    };

    unique case (NrLanes)
      1 : return lut_1lane [seqNbIdx][ew];
      2 : return lut_2lane [seqNbIdx][ew];
      4 : return lut_4lane [seqNbIdx][ew];
      8 : return lut_8lane [seqNbIdx][ew];
      16: return lut_16lane[seqNbIdx][ew];
      default: return 0;
	  endcase
  endfunction

  function automatic logic [{$clog2(riva_pkg::DLEN*riva_pkg::MaxNrLanes/4)}-1:0] query_seq_idx(input int NrLanes, input int shfNbIdx, input riscv_mv_pkg::vew_e ew);
    automatic logic [5-1:0] lut_1lane [0:31][0:3] = '{
      '{5'd000, 5'd000, 5'd000, 5'd000}, '{5'd016, 5'd001, 5'd001, 5'd001}, '{5'd008, 5'd016, 5'd002, 5'd002}, '{5'd024, 5'd017, 5'd003, 5'd003}, '{5'd004, 5'd008, 5'd016, 5'd004}, '{5'd020, 5'd009, 5'd017, 5'd005}, '{5'd012, 5'd024, 5'd018, 5'd006}, '{5'd028, 5'd025, 5'd019, 5'd007},
      '{5'd001, 5'd002, 5'd004, 5'd008}, '{5'd017, 5'd003, 5'd005, 5'd009}, '{5'd009, 5'd018, 5'd006, 5'd010}, '{5'd025, 5'd019, 5'd007, 5'd011}, '{5'd005, 5'd010, 5'd020, 5'd012}, '{5'd021, 5'd011, 5'd021, 5'd013}, '{5'd013, 5'd026, 5'd022, 5'd014}, '{5'd029, 5'd027, 5'd023, 5'd015},
      '{5'd002, 5'd004, 5'd008, 5'd016}, '{5'd018, 5'd005, 5'd009, 5'd017}, '{5'd010, 5'd020, 5'd010, 5'd018}, '{5'd026, 5'd021, 5'd011, 5'd019}, '{5'd006, 5'd012, 5'd024, 5'd020}, '{5'd022, 5'd013, 5'd025, 5'd021}, '{5'd014, 5'd028, 5'd026, 5'd022}, '{5'd030, 5'd029, 5'd027, 5'd023},
      '{5'd003, 5'd006, 5'd012, 5'd024}, '{5'd019, 5'd007, 5'd013, 5'd025}, '{5'd011, 5'd022, 5'd014, 5'd026}, '{5'd027, 5'd023, 5'd015, 5'd027}, '{5'd007, 5'd014, 5'd028, 5'd028}, '{5'd023, 5'd015, 5'd029, 5'd029}, '{5'd015, 5'd030, 5'd030, 5'd030}, '{5'd031, 5'd031, 5'd031, 5'd031}
    };
    automatic logic [6-1:0] lut_2lane [0:63][0:3] = '{
      '{6'd000, 6'd000, 6'd000, 6'd000}, '{6'd032, 6'd001, 6'd001, 6'd001}, '{6'd016, 6'd032, 6'd002, 6'd002}, '{6'd048, 6'd033, 6'd003, 6'd003}, '{6'd008, 6'd016, 6'd032, 6'd004}, '{6'd040, 6'd017, 6'd033, 6'd005}, '{6'd024, 6'd048, 6'd034, 6'd006}, '{6'd056, 6'd049, 6'd035, 6'd007},
      '{6'd002, 6'd004, 6'd008, 6'd016}, '{6'd034, 6'd005, 6'd009, 6'd017}, '{6'd018, 6'd036, 6'd010, 6'd018}, '{6'd050, 6'd037, 6'd011, 6'd019}, '{6'd010, 6'd020, 6'd040, 6'd020}, '{6'd042, 6'd021, 6'd041, 6'd021}, '{6'd026, 6'd052, 6'd042, 6'd022}, '{6'd058, 6'd053, 6'd043, 6'd023},
      '{6'd004, 6'd008, 6'd016, 6'd032}, '{6'd036, 6'd009, 6'd017, 6'd033}, '{6'd020, 6'd040, 6'd018, 6'd034}, '{6'd052, 6'd041, 6'd019, 6'd035}, '{6'd012, 6'd024, 6'd048, 6'd036}, '{6'd044, 6'd025, 6'd049, 6'd037}, '{6'd028, 6'd056, 6'd050, 6'd038}, '{6'd060, 6'd057, 6'd051, 6'd039},
      '{6'd006, 6'd012, 6'd024, 6'd048}, '{6'd038, 6'd013, 6'd025, 6'd049}, '{6'd022, 6'd044, 6'd026, 6'd050}, '{6'd054, 6'd045, 6'd027, 6'd051}, '{6'd014, 6'd028, 6'd056, 6'd052}, '{6'd046, 6'd029, 6'd057, 6'd053}, '{6'd030, 6'd060, 6'd058, 6'd054}, '{6'd062, 6'd061, 6'd059, 6'd055},
      '{6'd001, 6'd002, 6'd004, 6'd008}, '{6'd033, 6'd003, 6'd005, 6'd009}, '{6'd017, 6'd034, 6'd006, 6'd010}, '{6'd049, 6'd035, 6'd007, 6'd011}, '{6'd009, 6'd018, 6'd036, 6'd012}, '{6'd041, 6'd019, 6'd037, 6'd013}, '{6'd025, 6'd050, 6'd038, 6'd014}, '{6'd057, 6'd051, 6'd039, 6'd015},
      '{6'd003, 6'd006, 6'd012, 6'd024}, '{6'd035, 6'd007, 6'd013, 6'd025}, '{6'd019, 6'd038, 6'd014, 6'd026}, '{6'd051, 6'd039, 6'd015, 6'd027}, '{6'd011, 6'd022, 6'd044, 6'd028}, '{6'd043, 6'd023, 6'd045, 6'd029}, '{6'd027, 6'd054, 6'd046, 6'd030}, '{6'd059, 6'd055, 6'd047, 6'd031},
      '{6'd005, 6'd010, 6'd020, 6'd040}, '{6'd037, 6'd011, 6'd021, 6'd041}, '{6'd021, 6'd042, 6'd022, 6'd042}, '{6'd053, 6'd043, 6'd023, 6'd043}, '{6'd013, 6'd026, 6'd052, 6'd044}, '{6'd045, 6'd027, 6'd053, 6'd045}, '{6'd029, 6'd058, 6'd054, 6'd046}, '{6'd061, 6'd059, 6'd055, 6'd047},
      '{6'd007, 6'd014, 6'd028, 6'd056}, '{6'd039, 6'd015, 6'd029, 6'd057}, '{6'd023, 6'd046, 6'd030, 6'd058}, '{6'd055, 6'd047, 6'd031, 6'd059}, '{6'd015, 6'd030, 6'd060, 6'd060}, '{6'd047, 6'd031, 6'd061, 6'd061}, '{6'd031, 6'd062, 6'd062, 6'd062}, '{6'd063, 6'd063, 6'd063, 6'd063}
    };
    automatic logic [7-1:0] lut_4lane [0:127][0:3] = '{
      '{7'd000, 7'd000, 7'd000, 7'd000}, '{7'd064, 7'd001, 7'd001, 7'd001}, '{7'd032, 7'd064, 7'd002, 7'd002}, '{7'd096, 7'd065, 7'd003, 7'd003}, '{7'd016, 7'd032, 7'd064, 7'd004}, '{7'd080, 7'd033, 7'd065, 7'd005}, '{7'd048, 7'd096, 7'd066, 7'd006}, '{7'd112, 7'd097, 7'd067, 7'd007},
      '{7'd004, 7'd008, 7'd016, 7'd032}, '{7'd068, 7'd009, 7'd017, 7'd033}, '{7'd036, 7'd072, 7'd018, 7'd034}, '{7'd100, 7'd073, 7'd019, 7'd035}, '{7'd020, 7'd040, 7'd080, 7'd036}, '{7'd084, 7'd041, 7'd081, 7'd037}, '{7'd052, 7'd104, 7'd082, 7'd038}, '{7'd116, 7'd105, 7'd083, 7'd039},
      '{7'd008, 7'd016, 7'd032, 7'd064}, '{7'd072, 7'd017, 7'd033, 7'd065}, '{7'd040, 7'd080, 7'd034, 7'd066}, '{7'd104, 7'd081, 7'd035, 7'd067}, '{7'd024, 7'd048, 7'd096, 7'd068}, '{7'd088, 7'd049, 7'd097, 7'd069}, '{7'd056, 7'd112, 7'd098, 7'd070}, '{7'd120, 7'd113, 7'd099, 7'd071},
      '{7'd012, 7'd024, 7'd048, 7'd096}, '{7'd076, 7'd025, 7'd049, 7'd097}, '{7'd044, 7'd088, 7'd050, 7'd098}, '{7'd108, 7'd089, 7'd051, 7'd099}, '{7'd028, 7'd056, 7'd112, 7'd100}, '{7'd092, 7'd057, 7'd113, 7'd101}, '{7'd060, 7'd120, 7'd114, 7'd102}, '{7'd124, 7'd121, 7'd115, 7'd103},
      '{7'd001, 7'd002, 7'd004, 7'd008}, '{7'd065, 7'd003, 7'd005, 7'd009}, '{7'd033, 7'd066, 7'd006, 7'd010}, '{7'd097, 7'd067, 7'd007, 7'd011}, '{7'd017, 7'd034, 7'd068, 7'd012}, '{7'd081, 7'd035, 7'd069, 7'd013}, '{7'd049, 7'd098, 7'd070, 7'd014}, '{7'd113, 7'd099, 7'd071, 7'd015},
      '{7'd005, 7'd010, 7'd020, 7'd040}, '{7'd069, 7'd011, 7'd021, 7'd041}, '{7'd037, 7'd074, 7'd022, 7'd042}, '{7'd101, 7'd075, 7'd023, 7'd043}, '{7'd021, 7'd042, 7'd084, 7'd044}, '{7'd085, 7'd043, 7'd085, 7'd045}, '{7'd053, 7'd106, 7'd086, 7'd046}, '{7'd117, 7'd107, 7'd087, 7'd047},
      '{7'd009, 7'd018, 7'd036, 7'd072}, '{7'd073, 7'd019, 7'd037, 7'd073}, '{7'd041, 7'd082, 7'd038, 7'd074}, '{7'd105, 7'd083, 7'd039, 7'd075}, '{7'd025, 7'd050, 7'd100, 7'd076}, '{7'd089, 7'd051, 7'd101, 7'd077}, '{7'd057, 7'd114, 7'd102, 7'd078}, '{7'd121, 7'd115, 7'd103, 7'd079},
      '{7'd013, 7'd026, 7'd052, 7'd104}, '{7'd077, 7'd027, 7'd053, 7'd105}, '{7'd045, 7'd090, 7'd054, 7'd106}, '{7'd109, 7'd091, 7'd055, 7'd107}, '{7'd029, 7'd058, 7'd116, 7'd108}, '{7'd093, 7'd059, 7'd117, 7'd109}, '{7'd061, 7'd122, 7'd118, 7'd110}, '{7'd125, 7'd123, 7'd119, 7'd111},
      '{7'd002, 7'd004, 7'd008, 7'd016}, '{7'd066, 7'd005, 7'd009, 7'd017}, '{7'd034, 7'd068, 7'd010, 7'd018}, '{7'd098, 7'd069, 7'd011, 7'd019}, '{7'd018, 7'd036, 7'd072, 7'd020}, '{7'd082, 7'd037, 7'd073, 7'd021}, '{7'd050, 7'd100, 7'd074, 7'd022}, '{7'd114, 7'd101, 7'd075, 7'd023},
      '{7'd006, 7'd012, 7'd024, 7'd048}, '{7'd070, 7'd013, 7'd025, 7'd049}, '{7'd038, 7'd076, 7'd026, 7'd050}, '{7'd102, 7'd077, 7'd027, 7'd051}, '{7'd022, 7'd044, 7'd088, 7'd052}, '{7'd086, 7'd045, 7'd089, 7'd053}, '{7'd054, 7'd108, 7'd090, 7'd054}, '{7'd118, 7'd109, 7'd091, 7'd055},
      '{7'd010, 7'd020, 7'd040, 7'd080}, '{7'd074, 7'd021, 7'd041, 7'd081}, '{7'd042, 7'd084, 7'd042, 7'd082}, '{7'd106, 7'd085, 7'd043, 7'd083}, '{7'd026, 7'd052, 7'd104, 7'd084}, '{7'd090, 7'd053, 7'd105, 7'd085}, '{7'd058, 7'd116, 7'd106, 7'd086}, '{7'd122, 7'd117, 7'd107, 7'd087},
      '{7'd014, 7'd028, 7'd056, 7'd112}, '{7'd078, 7'd029, 7'd057, 7'd113}, '{7'd046, 7'd092, 7'd058, 7'd114}, '{7'd110, 7'd093, 7'd059, 7'd115}, '{7'd030, 7'd060, 7'd120, 7'd116}, '{7'd094, 7'd061, 7'd121, 7'd117}, '{7'd062, 7'd124, 7'd122, 7'd118}, '{7'd126, 7'd125, 7'd123, 7'd119},
      '{7'd003, 7'd006, 7'd012, 7'd024}, '{7'd067, 7'd007, 7'd013, 7'd025}, '{7'd035, 7'd070, 7'd014, 7'd026}, '{7'd099, 7'd071, 7'd015, 7'd027}, '{7'd019, 7'd038, 7'd076, 7'd028}, '{7'd083, 7'd039, 7'd077, 7'd029}, '{7'd051, 7'd102, 7'd078, 7'd030}, '{7'd115, 7'd103, 7'd079, 7'd031},
      '{7'd007, 7'd014, 7'd028, 7'd056}, '{7'd071, 7'd015, 7'd029, 7'd057}, '{7'd039, 7'd078, 7'd030, 7'd058}, '{7'd103, 7'd079, 7'd031, 7'd059}, '{7'd023, 7'd046, 7'd092, 7'd060}, '{7'd087, 7'd047, 7'd093, 7'd061}, '{7'd055, 7'd110, 7'd094, 7'd062}, '{7'd119, 7'd111, 7'd095, 7'd063},
      '{7'd011, 7'd022, 7'd044, 7'd088}, '{7'd075, 7'd023, 7'd045, 7'd089}, '{7'd043, 7'd086, 7'd046, 7'd090}, '{7'd107, 7'd087, 7'd047, 7'd091}, '{7'd027, 7'd054, 7'd108, 7'd092}, '{7'd091, 7'd055, 7'd109, 7'd093}, '{7'd059, 7'd118, 7'd110, 7'd094}, '{7'd123, 7'd119, 7'd111, 7'd095},
      '{7'd015, 7'd030, 7'd060, 7'd120}, '{7'd079, 7'd031, 7'd061, 7'd121}, '{7'd047, 7'd094, 7'd062, 7'd122}, '{7'd111, 7'd095, 7'd063, 7'd123}, '{7'd031, 7'd062, 7'd124, 7'd124}, '{7'd095, 7'd063, 7'd125, 7'd125}, '{7'd063, 7'd126, 7'd126, 7'd126}, '{7'd127, 7'd127, 7'd127, 7'd127}
    };
    automatic logic [8-1:0] lut_8lane [0:255][0:3] = '{
      '{8'd000, 8'd000, 8'd000, 8'd000}, '{8'd128, 8'd001, 8'd001, 8'd001}, '{8'd064, 8'd128, 8'd002, 8'd002}, '{8'd192, 8'd129, 8'd003, 8'd003}, '{8'd032, 8'd064, 8'd128, 8'd004}, '{8'd160, 8'd065, 8'd129, 8'd005}, '{8'd096, 8'd192, 8'd130, 8'd006}, '{8'd224, 8'd193, 8'd131, 8'd007},
      '{8'd008, 8'd016, 8'd032, 8'd064}, '{8'd136, 8'd017, 8'd033, 8'd065}, '{8'd072, 8'd144, 8'd034, 8'd066}, '{8'd200, 8'd145, 8'd035, 8'd067}, '{8'd040, 8'd080, 8'd160, 8'd068}, '{8'd168, 8'd081, 8'd161, 8'd069}, '{8'd104, 8'd208, 8'd162, 8'd070}, '{8'd232, 8'd209, 8'd163, 8'd071},
      '{8'd016, 8'd032, 8'd064, 8'd128}, '{8'd144, 8'd033, 8'd065, 8'd129}, '{8'd080, 8'd160, 8'd066, 8'd130}, '{8'd208, 8'd161, 8'd067, 8'd131}, '{8'd048, 8'd096, 8'd192, 8'd132}, '{8'd176, 8'd097, 8'd193, 8'd133}, '{8'd112, 8'd224, 8'd194, 8'd134}, '{8'd240, 8'd225, 8'd195, 8'd135},
      '{8'd024, 8'd048, 8'd096, 8'd192}, '{8'd152, 8'd049, 8'd097, 8'd193}, '{8'd088, 8'd176, 8'd098, 8'd194}, '{8'd216, 8'd177, 8'd099, 8'd195}, '{8'd056, 8'd112, 8'd224, 8'd196}, '{8'd184, 8'd113, 8'd225, 8'd197}, '{8'd120, 8'd240, 8'd226, 8'd198}, '{8'd248, 8'd241, 8'd227, 8'd199},
      '{8'd001, 8'd002, 8'd004, 8'd008}, '{8'd129, 8'd003, 8'd005, 8'd009}, '{8'd065, 8'd130, 8'd006, 8'd010}, '{8'd193, 8'd131, 8'd007, 8'd011}, '{8'd033, 8'd066, 8'd132, 8'd012}, '{8'd161, 8'd067, 8'd133, 8'd013}, '{8'd097, 8'd194, 8'd134, 8'd014}, '{8'd225, 8'd195, 8'd135, 8'd015},
      '{8'd009, 8'd018, 8'd036, 8'd072}, '{8'd137, 8'd019, 8'd037, 8'd073}, '{8'd073, 8'd146, 8'd038, 8'd074}, '{8'd201, 8'd147, 8'd039, 8'd075}, '{8'd041, 8'd082, 8'd164, 8'd076}, '{8'd169, 8'd083, 8'd165, 8'd077}, '{8'd105, 8'd210, 8'd166, 8'd078}, '{8'd233, 8'd211, 8'd167, 8'd079},
      '{8'd017, 8'd034, 8'd068, 8'd136}, '{8'd145, 8'd035, 8'd069, 8'd137}, '{8'd081, 8'd162, 8'd070, 8'd138}, '{8'd209, 8'd163, 8'd071, 8'd139}, '{8'd049, 8'd098, 8'd196, 8'd140}, '{8'd177, 8'd099, 8'd197, 8'd141}, '{8'd113, 8'd226, 8'd198, 8'd142}, '{8'd241, 8'd227, 8'd199, 8'd143},
      '{8'd025, 8'd050, 8'd100, 8'd200}, '{8'd153, 8'd051, 8'd101, 8'd201}, '{8'd089, 8'd178, 8'd102, 8'd202}, '{8'd217, 8'd179, 8'd103, 8'd203}, '{8'd057, 8'd114, 8'd228, 8'd204}, '{8'd185, 8'd115, 8'd229, 8'd205}, '{8'd121, 8'd242, 8'd230, 8'd206}, '{8'd249, 8'd243, 8'd231, 8'd207},
      '{8'd002, 8'd004, 8'd008, 8'd016}, '{8'd130, 8'd005, 8'd009, 8'd017}, '{8'd066, 8'd132, 8'd010, 8'd018}, '{8'd194, 8'd133, 8'd011, 8'd019}, '{8'd034, 8'd068, 8'd136, 8'd020}, '{8'd162, 8'd069, 8'd137, 8'd021}, '{8'd098, 8'd196, 8'd138, 8'd022}, '{8'd226, 8'd197, 8'd139, 8'd023},
      '{8'd010, 8'd020, 8'd040, 8'd080}, '{8'd138, 8'd021, 8'd041, 8'd081}, '{8'd074, 8'd148, 8'd042, 8'd082}, '{8'd202, 8'd149, 8'd043, 8'd083}, '{8'd042, 8'd084, 8'd168, 8'd084}, '{8'd170, 8'd085, 8'd169, 8'd085}, '{8'd106, 8'd212, 8'd170, 8'd086}, '{8'd234, 8'd213, 8'd171, 8'd087},
      '{8'd018, 8'd036, 8'd072, 8'd144}, '{8'd146, 8'd037, 8'd073, 8'd145}, '{8'd082, 8'd164, 8'd074, 8'd146}, '{8'd210, 8'd165, 8'd075, 8'd147}, '{8'd050, 8'd100, 8'd200, 8'd148}, '{8'd178, 8'd101, 8'd201, 8'd149}, '{8'd114, 8'd228, 8'd202, 8'd150}, '{8'd242, 8'd229, 8'd203, 8'd151},
      '{8'd026, 8'd052, 8'd104, 8'd208}, '{8'd154, 8'd053, 8'd105, 8'd209}, '{8'd090, 8'd180, 8'd106, 8'd210}, '{8'd218, 8'd181, 8'd107, 8'd211}, '{8'd058, 8'd116, 8'd232, 8'd212}, '{8'd186, 8'd117, 8'd233, 8'd213}, '{8'd122, 8'd244, 8'd234, 8'd214}, '{8'd250, 8'd245, 8'd235, 8'd215},
      '{8'd003, 8'd006, 8'd012, 8'd024}, '{8'd131, 8'd007, 8'd013, 8'd025}, '{8'd067, 8'd134, 8'd014, 8'd026}, '{8'd195, 8'd135, 8'd015, 8'd027}, '{8'd035, 8'd070, 8'd140, 8'd028}, '{8'd163, 8'd071, 8'd141, 8'd029}, '{8'd099, 8'd198, 8'd142, 8'd030}, '{8'd227, 8'd199, 8'd143, 8'd031},
      '{8'd011, 8'd022, 8'd044, 8'd088}, '{8'd139, 8'd023, 8'd045, 8'd089}, '{8'd075, 8'd150, 8'd046, 8'd090}, '{8'd203, 8'd151, 8'd047, 8'd091}, '{8'd043, 8'd086, 8'd172, 8'd092}, '{8'd171, 8'd087, 8'd173, 8'd093}, '{8'd107, 8'd214, 8'd174, 8'd094}, '{8'd235, 8'd215, 8'd175, 8'd095},
      '{8'd019, 8'd038, 8'd076, 8'd152}, '{8'd147, 8'd039, 8'd077, 8'd153}, '{8'd083, 8'd166, 8'd078, 8'd154}, '{8'd211, 8'd167, 8'd079, 8'd155}, '{8'd051, 8'd102, 8'd204, 8'd156}, '{8'd179, 8'd103, 8'd205, 8'd157}, '{8'd115, 8'd230, 8'd206, 8'd158}, '{8'd243, 8'd231, 8'd207, 8'd159},
      '{8'd027, 8'd054, 8'd108, 8'd216}, '{8'd155, 8'd055, 8'd109, 8'd217}, '{8'd091, 8'd182, 8'd110, 8'd218}, '{8'd219, 8'd183, 8'd111, 8'd219}, '{8'd059, 8'd118, 8'd236, 8'd220}, '{8'd187, 8'd119, 8'd237, 8'd221}, '{8'd123, 8'd246, 8'd238, 8'd222}, '{8'd251, 8'd247, 8'd239, 8'd223},
      '{8'd004, 8'd008, 8'd016, 8'd032}, '{8'd132, 8'd009, 8'd017, 8'd033}, '{8'd068, 8'd136, 8'd018, 8'd034}, '{8'd196, 8'd137, 8'd019, 8'd035}, '{8'd036, 8'd072, 8'd144, 8'd036}, '{8'd164, 8'd073, 8'd145, 8'd037}, '{8'd100, 8'd200, 8'd146, 8'd038}, '{8'd228, 8'd201, 8'd147, 8'd039},
      '{8'd012, 8'd024, 8'd048, 8'd096}, '{8'd140, 8'd025, 8'd049, 8'd097}, '{8'd076, 8'd152, 8'd050, 8'd098}, '{8'd204, 8'd153, 8'd051, 8'd099}, '{8'd044, 8'd088, 8'd176, 8'd100}, '{8'd172, 8'd089, 8'd177, 8'd101}, '{8'd108, 8'd216, 8'd178, 8'd102}, '{8'd236, 8'd217, 8'd179, 8'd103},
      '{8'd020, 8'd040, 8'd080, 8'd160}, '{8'd148, 8'd041, 8'd081, 8'd161}, '{8'd084, 8'd168, 8'd082, 8'd162}, '{8'd212, 8'd169, 8'd083, 8'd163}, '{8'd052, 8'd104, 8'd208, 8'd164}, '{8'd180, 8'd105, 8'd209, 8'd165}, '{8'd116, 8'd232, 8'd210, 8'd166}, '{8'd244, 8'd233, 8'd211, 8'd167},
      '{8'd028, 8'd056, 8'd112, 8'd224}, '{8'd156, 8'd057, 8'd113, 8'd225}, '{8'd092, 8'd184, 8'd114, 8'd226}, '{8'd220, 8'd185, 8'd115, 8'd227}, '{8'd060, 8'd120, 8'd240, 8'd228}, '{8'd188, 8'd121, 8'd241, 8'd229}, '{8'd124, 8'd248, 8'd242, 8'd230}, '{8'd252, 8'd249, 8'd243, 8'd231},
      '{8'd005, 8'd010, 8'd020, 8'd040}, '{8'd133, 8'd011, 8'd021, 8'd041}, '{8'd069, 8'd138, 8'd022, 8'd042}, '{8'd197, 8'd139, 8'd023, 8'd043}, '{8'd037, 8'd074, 8'd148, 8'd044}, '{8'd165, 8'd075, 8'd149, 8'd045}, '{8'd101, 8'd202, 8'd150, 8'd046}, '{8'd229, 8'd203, 8'd151, 8'd047},
      '{8'd013, 8'd026, 8'd052, 8'd104}, '{8'd141, 8'd027, 8'd053, 8'd105}, '{8'd077, 8'd154, 8'd054, 8'd106}, '{8'd205, 8'd155, 8'd055, 8'd107}, '{8'd045, 8'd090, 8'd180, 8'd108}, '{8'd173, 8'd091, 8'd181, 8'd109}, '{8'd109, 8'd218, 8'd182, 8'd110}, '{8'd237, 8'd219, 8'd183, 8'd111},
      '{8'd021, 8'd042, 8'd084, 8'd168}, '{8'd149, 8'd043, 8'd085, 8'd169}, '{8'd085, 8'd170, 8'd086, 8'd170}, '{8'd213, 8'd171, 8'd087, 8'd171}, '{8'd053, 8'd106, 8'd212, 8'd172}, '{8'd181, 8'd107, 8'd213, 8'd173}, '{8'd117, 8'd234, 8'd214, 8'd174}, '{8'd245, 8'd235, 8'd215, 8'd175},
      '{8'd029, 8'd058, 8'd116, 8'd232}, '{8'd157, 8'd059, 8'd117, 8'd233}, '{8'd093, 8'd186, 8'd118, 8'd234}, '{8'd221, 8'd187, 8'd119, 8'd235}, '{8'd061, 8'd122, 8'd244, 8'd236}, '{8'd189, 8'd123, 8'd245, 8'd237}, '{8'd125, 8'd250, 8'd246, 8'd238}, '{8'd253, 8'd251, 8'd247, 8'd239},
      '{8'd006, 8'd012, 8'd024, 8'd048}, '{8'd134, 8'd013, 8'd025, 8'd049}, '{8'd070, 8'd140, 8'd026, 8'd050}, '{8'd198, 8'd141, 8'd027, 8'd051}, '{8'd038, 8'd076, 8'd152, 8'd052}, '{8'd166, 8'd077, 8'd153, 8'd053}, '{8'd102, 8'd204, 8'd154, 8'd054}, '{8'd230, 8'd205, 8'd155, 8'd055},
      '{8'd014, 8'd028, 8'd056, 8'd112}, '{8'd142, 8'd029, 8'd057, 8'd113}, '{8'd078, 8'd156, 8'd058, 8'd114}, '{8'd206, 8'd157, 8'd059, 8'd115}, '{8'd046, 8'd092, 8'd184, 8'd116}, '{8'd174, 8'd093, 8'd185, 8'd117}, '{8'd110, 8'd220, 8'd186, 8'd118}, '{8'd238, 8'd221, 8'd187, 8'd119},
      '{8'd022, 8'd044, 8'd088, 8'd176}, '{8'd150, 8'd045, 8'd089, 8'd177}, '{8'd086, 8'd172, 8'd090, 8'd178}, '{8'd214, 8'd173, 8'd091, 8'd179}, '{8'd054, 8'd108, 8'd216, 8'd180}, '{8'd182, 8'd109, 8'd217, 8'd181}, '{8'd118, 8'd236, 8'd218, 8'd182}, '{8'd246, 8'd237, 8'd219, 8'd183},
      '{8'd030, 8'd060, 8'd120, 8'd240}, '{8'd158, 8'd061, 8'd121, 8'd241}, '{8'd094, 8'd188, 8'd122, 8'd242}, '{8'd222, 8'd189, 8'd123, 8'd243}, '{8'd062, 8'd124, 8'd248, 8'd244}, '{8'd190, 8'd125, 8'd249, 8'd245}, '{8'd126, 8'd252, 8'd250, 8'd246}, '{8'd254, 8'd253, 8'd251, 8'd247},
      '{8'd007, 8'd014, 8'd028, 8'd056}, '{8'd135, 8'd015, 8'd029, 8'd057}, '{8'd071, 8'd142, 8'd030, 8'd058}, '{8'd199, 8'd143, 8'd031, 8'd059}, '{8'd039, 8'd078, 8'd156, 8'd060}, '{8'd167, 8'd079, 8'd157, 8'd061}, '{8'd103, 8'd206, 8'd158, 8'd062}, '{8'd231, 8'd207, 8'd159, 8'd063},
      '{8'd015, 8'd030, 8'd060, 8'd120}, '{8'd143, 8'd031, 8'd061, 8'd121}, '{8'd079, 8'd158, 8'd062, 8'd122}, '{8'd207, 8'd159, 8'd063, 8'd123}, '{8'd047, 8'd094, 8'd188, 8'd124}, '{8'd175, 8'd095, 8'd189, 8'd125}, '{8'd111, 8'd222, 8'd190, 8'd126}, '{8'd239, 8'd223, 8'd191, 8'd127},
      '{8'd023, 8'd046, 8'd092, 8'd184}, '{8'd151, 8'd047, 8'd093, 8'd185}, '{8'd087, 8'd174, 8'd094, 8'd186}, '{8'd215, 8'd175, 8'd095, 8'd187}, '{8'd055, 8'd110, 8'd220, 8'd188}, '{8'd183, 8'd111, 8'd221, 8'd189}, '{8'd119, 8'd238, 8'd222, 8'd190}, '{8'd247, 8'd239, 8'd223, 8'd191},
      '{8'd031, 8'd062, 8'd124, 8'd248}, '{8'd159, 8'd063, 8'd125, 8'd249}, '{8'd095, 8'd190, 8'd126, 8'd250}, '{8'd223, 8'd191, 8'd127, 8'd251}, '{8'd063, 8'd126, 8'd252, 8'd252}, '{8'd191, 8'd127, 8'd253, 8'd253}, '{8'd127, 8'd254, 8'd254, 8'd254}, '{8'd255, 8'd255, 8'd255, 8'd255}
    };
    automatic logic [9-1:0] lut_16lane [0:511][0:3] = '{
      '{9'd000, 9'd000, 9'd000, 9'd000}, '{9'd256, 9'd001, 9'd001, 9'd001}, '{9'd128, 9'd256, 9'd002, 9'd002}, '{9'd384, 9'd257, 9'd003, 9'd003}, '{9'd064, 9'd128, 9'd256, 9'd004}, '{9'd320, 9'd129, 9'd257, 9'd005}, '{9'd192, 9'd384, 9'd258, 9'd006}, '{9'd448, 9'd385, 9'd259, 9'd007},
      '{9'd016, 9'd032, 9'd064, 9'd128}, '{9'd272, 9'd033, 9'd065, 9'd129}, '{9'd144, 9'd288, 9'd066, 9'd130}, '{9'd400, 9'd289, 9'd067, 9'd131}, '{9'd080, 9'd160, 9'd320, 9'd132}, '{9'd336, 9'd161, 9'd321, 9'd133}, '{9'd208, 9'd416, 9'd322, 9'd134}, '{9'd464, 9'd417, 9'd323, 9'd135},
      '{9'd032, 9'd064, 9'd128, 9'd256}, '{9'd288, 9'd065, 9'd129, 9'd257}, '{9'd160, 9'd320, 9'd130, 9'd258}, '{9'd416, 9'd321, 9'd131, 9'd259}, '{9'd096, 9'd192, 9'd384, 9'd260}, '{9'd352, 9'd193, 9'd385, 9'd261}, '{9'd224, 9'd448, 9'd386, 9'd262}, '{9'd480, 9'd449, 9'd387, 9'd263},
      '{9'd048, 9'd096, 9'd192, 9'd384}, '{9'd304, 9'd097, 9'd193, 9'd385}, '{9'd176, 9'd352, 9'd194, 9'd386}, '{9'd432, 9'd353, 9'd195, 9'd387}, '{9'd112, 9'd224, 9'd448, 9'd388}, '{9'd368, 9'd225, 9'd449, 9'd389}, '{9'd240, 9'd480, 9'd450, 9'd390}, '{9'd496, 9'd481, 9'd451, 9'd391},
      '{9'd001, 9'd002, 9'd004, 9'd008}, '{9'd257, 9'd003, 9'd005, 9'd009}, '{9'd129, 9'd258, 9'd006, 9'd010}, '{9'd385, 9'd259, 9'd007, 9'd011}, '{9'd065, 9'd130, 9'd260, 9'd012}, '{9'd321, 9'd131, 9'd261, 9'd013}, '{9'd193, 9'd386, 9'd262, 9'd014}, '{9'd449, 9'd387, 9'd263, 9'd015},
      '{9'd017, 9'd034, 9'd068, 9'd136}, '{9'd273, 9'd035, 9'd069, 9'd137}, '{9'd145, 9'd290, 9'd070, 9'd138}, '{9'd401, 9'd291, 9'd071, 9'd139}, '{9'd081, 9'd162, 9'd324, 9'd140}, '{9'd337, 9'd163, 9'd325, 9'd141}, '{9'd209, 9'd418, 9'd326, 9'd142}, '{9'd465, 9'd419, 9'd327, 9'd143},
      '{9'd033, 9'd066, 9'd132, 9'd264}, '{9'd289, 9'd067, 9'd133, 9'd265}, '{9'd161, 9'd322, 9'd134, 9'd266}, '{9'd417, 9'd323, 9'd135, 9'd267}, '{9'd097, 9'd194, 9'd388, 9'd268}, '{9'd353, 9'd195, 9'd389, 9'd269}, '{9'd225, 9'd450, 9'd390, 9'd270}, '{9'd481, 9'd451, 9'd391, 9'd271},
      '{9'd049, 9'd098, 9'd196, 9'd392}, '{9'd305, 9'd099, 9'd197, 9'd393}, '{9'd177, 9'd354, 9'd198, 9'd394}, '{9'd433, 9'd355, 9'd199, 9'd395}, '{9'd113, 9'd226, 9'd452, 9'd396}, '{9'd369, 9'd227, 9'd453, 9'd397}, '{9'd241, 9'd482, 9'd454, 9'd398}, '{9'd497, 9'd483, 9'd455, 9'd399},
      '{9'd002, 9'd004, 9'd008, 9'd016}, '{9'd258, 9'd005, 9'd009, 9'd017}, '{9'd130, 9'd260, 9'd010, 9'd018}, '{9'd386, 9'd261, 9'd011, 9'd019}, '{9'd066, 9'd132, 9'd264, 9'd020}, '{9'd322, 9'd133, 9'd265, 9'd021}, '{9'd194, 9'd388, 9'd266, 9'd022}, '{9'd450, 9'd389, 9'd267, 9'd023},
      '{9'd018, 9'd036, 9'd072, 9'd144}, '{9'd274, 9'd037, 9'd073, 9'd145}, '{9'd146, 9'd292, 9'd074, 9'd146}, '{9'd402, 9'd293, 9'd075, 9'd147}, '{9'd082, 9'd164, 9'd328, 9'd148}, '{9'd338, 9'd165, 9'd329, 9'd149}, '{9'd210, 9'd420, 9'd330, 9'd150}, '{9'd466, 9'd421, 9'd331, 9'd151},
      '{9'd034, 9'd068, 9'd136, 9'd272}, '{9'd290, 9'd069, 9'd137, 9'd273}, '{9'd162, 9'd324, 9'd138, 9'd274}, '{9'd418, 9'd325, 9'd139, 9'd275}, '{9'd098, 9'd196, 9'd392, 9'd276}, '{9'd354, 9'd197, 9'd393, 9'd277}, '{9'd226, 9'd452, 9'd394, 9'd278}, '{9'd482, 9'd453, 9'd395, 9'd279},
      '{9'd050, 9'd100, 9'd200, 9'd400}, '{9'd306, 9'd101, 9'd201, 9'd401}, '{9'd178, 9'd356, 9'd202, 9'd402}, '{9'd434, 9'd357, 9'd203, 9'd403}, '{9'd114, 9'd228, 9'd456, 9'd404}, '{9'd370, 9'd229, 9'd457, 9'd405}, '{9'd242, 9'd484, 9'd458, 9'd406}, '{9'd498, 9'd485, 9'd459, 9'd407},
      '{9'd003, 9'd006, 9'd012, 9'd024}, '{9'd259, 9'd007, 9'd013, 9'd025}, '{9'd131, 9'd262, 9'd014, 9'd026}, '{9'd387, 9'd263, 9'd015, 9'd027}, '{9'd067, 9'd134, 9'd268, 9'd028}, '{9'd323, 9'd135, 9'd269, 9'd029}, '{9'd195, 9'd390, 9'd270, 9'd030}, '{9'd451, 9'd391, 9'd271, 9'd031},
      '{9'd019, 9'd038, 9'd076, 9'd152}, '{9'd275, 9'd039, 9'd077, 9'd153}, '{9'd147, 9'd294, 9'd078, 9'd154}, '{9'd403, 9'd295, 9'd079, 9'd155}, '{9'd083, 9'd166, 9'd332, 9'd156}, '{9'd339, 9'd167, 9'd333, 9'd157}, '{9'd211, 9'd422, 9'd334, 9'd158}, '{9'd467, 9'd423, 9'd335, 9'd159},
      '{9'd035, 9'd070, 9'd140, 9'd280}, '{9'd291, 9'd071, 9'd141, 9'd281}, '{9'd163, 9'd326, 9'd142, 9'd282}, '{9'd419, 9'd327, 9'd143, 9'd283}, '{9'd099, 9'd198, 9'd396, 9'd284}, '{9'd355, 9'd199, 9'd397, 9'd285}, '{9'd227, 9'd454, 9'd398, 9'd286}, '{9'd483, 9'd455, 9'd399, 9'd287},
      '{9'd051, 9'd102, 9'd204, 9'd408}, '{9'd307, 9'd103, 9'd205, 9'd409}, '{9'd179, 9'd358, 9'd206, 9'd410}, '{9'd435, 9'd359, 9'd207, 9'd411}, '{9'd115, 9'd230, 9'd460, 9'd412}, '{9'd371, 9'd231, 9'd461, 9'd413}, '{9'd243, 9'd486, 9'd462, 9'd414}, '{9'd499, 9'd487, 9'd463, 9'd415},
      '{9'd004, 9'd008, 9'd016, 9'd032}, '{9'd260, 9'd009, 9'd017, 9'd033}, '{9'd132, 9'd264, 9'd018, 9'd034}, '{9'd388, 9'd265, 9'd019, 9'd035}, '{9'd068, 9'd136, 9'd272, 9'd036}, '{9'd324, 9'd137, 9'd273, 9'd037}, '{9'd196, 9'd392, 9'd274, 9'd038}, '{9'd452, 9'd393, 9'd275, 9'd039},
      '{9'd020, 9'd040, 9'd080, 9'd160}, '{9'd276, 9'd041, 9'd081, 9'd161}, '{9'd148, 9'd296, 9'd082, 9'd162}, '{9'd404, 9'd297, 9'd083, 9'd163}, '{9'd084, 9'd168, 9'd336, 9'd164}, '{9'd340, 9'd169, 9'd337, 9'd165}, '{9'd212, 9'd424, 9'd338, 9'd166}, '{9'd468, 9'd425, 9'd339, 9'd167},
      '{9'd036, 9'd072, 9'd144, 9'd288}, '{9'd292, 9'd073, 9'd145, 9'd289}, '{9'd164, 9'd328, 9'd146, 9'd290}, '{9'd420, 9'd329, 9'd147, 9'd291}, '{9'd100, 9'd200, 9'd400, 9'd292}, '{9'd356, 9'd201, 9'd401, 9'd293}, '{9'd228, 9'd456, 9'd402, 9'd294}, '{9'd484, 9'd457, 9'd403, 9'd295},
      '{9'd052, 9'd104, 9'd208, 9'd416}, '{9'd308, 9'd105, 9'd209, 9'd417}, '{9'd180, 9'd360, 9'd210, 9'd418}, '{9'd436, 9'd361, 9'd211, 9'd419}, '{9'd116, 9'd232, 9'd464, 9'd420}, '{9'd372, 9'd233, 9'd465, 9'd421}, '{9'd244, 9'd488, 9'd466, 9'd422}, '{9'd500, 9'd489, 9'd467, 9'd423},
      '{9'd005, 9'd010, 9'd020, 9'd040}, '{9'd261, 9'd011, 9'd021, 9'd041}, '{9'd133, 9'd266, 9'd022, 9'd042}, '{9'd389, 9'd267, 9'd023, 9'd043}, '{9'd069, 9'd138, 9'd276, 9'd044}, '{9'd325, 9'd139, 9'd277, 9'd045}, '{9'd197, 9'd394, 9'd278, 9'd046}, '{9'd453, 9'd395, 9'd279, 9'd047},
      '{9'd021, 9'd042, 9'd084, 9'd168}, '{9'd277, 9'd043, 9'd085, 9'd169}, '{9'd149, 9'd298, 9'd086, 9'd170}, '{9'd405, 9'd299, 9'd087, 9'd171}, '{9'd085, 9'd170, 9'd340, 9'd172}, '{9'd341, 9'd171, 9'd341, 9'd173}, '{9'd213, 9'd426, 9'd342, 9'd174}, '{9'd469, 9'd427, 9'd343, 9'd175},
      '{9'd037, 9'd074, 9'd148, 9'd296}, '{9'd293, 9'd075, 9'd149, 9'd297}, '{9'd165, 9'd330, 9'd150, 9'd298}, '{9'd421, 9'd331, 9'd151, 9'd299}, '{9'd101, 9'd202, 9'd404, 9'd300}, '{9'd357, 9'd203, 9'd405, 9'd301}, '{9'd229, 9'd458, 9'd406, 9'd302}, '{9'd485, 9'd459, 9'd407, 9'd303},
      '{9'd053, 9'd106, 9'd212, 9'd424}, '{9'd309, 9'd107, 9'd213, 9'd425}, '{9'd181, 9'd362, 9'd214, 9'd426}, '{9'd437, 9'd363, 9'd215, 9'd427}, '{9'd117, 9'd234, 9'd468, 9'd428}, '{9'd373, 9'd235, 9'd469, 9'd429}, '{9'd245, 9'd490, 9'd470, 9'd430}, '{9'd501, 9'd491, 9'd471, 9'd431},
      '{9'd006, 9'd012, 9'd024, 9'd048}, '{9'd262, 9'd013, 9'd025, 9'd049}, '{9'd134, 9'd268, 9'd026, 9'd050}, '{9'd390, 9'd269, 9'd027, 9'd051}, '{9'd070, 9'd140, 9'd280, 9'd052}, '{9'd326, 9'd141, 9'd281, 9'd053}, '{9'd198, 9'd396, 9'd282, 9'd054}, '{9'd454, 9'd397, 9'd283, 9'd055},
      '{9'd022, 9'd044, 9'd088, 9'd176}, '{9'd278, 9'd045, 9'd089, 9'd177}, '{9'd150, 9'd300, 9'd090, 9'd178}, '{9'd406, 9'd301, 9'd091, 9'd179}, '{9'd086, 9'd172, 9'd344, 9'd180}, '{9'd342, 9'd173, 9'd345, 9'd181}, '{9'd214, 9'd428, 9'd346, 9'd182}, '{9'd470, 9'd429, 9'd347, 9'd183},
      '{9'd038, 9'd076, 9'd152, 9'd304}, '{9'd294, 9'd077, 9'd153, 9'd305}, '{9'd166, 9'd332, 9'd154, 9'd306}, '{9'd422, 9'd333, 9'd155, 9'd307}, '{9'd102, 9'd204, 9'd408, 9'd308}, '{9'd358, 9'd205, 9'd409, 9'd309}, '{9'd230, 9'd460, 9'd410, 9'd310}, '{9'd486, 9'd461, 9'd411, 9'd311},
      '{9'd054, 9'd108, 9'd216, 9'd432}, '{9'd310, 9'd109, 9'd217, 9'd433}, '{9'd182, 9'd364, 9'd218, 9'd434}, '{9'd438, 9'd365, 9'd219, 9'd435}, '{9'd118, 9'd236, 9'd472, 9'd436}, '{9'd374, 9'd237, 9'd473, 9'd437}, '{9'd246, 9'd492, 9'd474, 9'd438}, '{9'd502, 9'd493, 9'd475, 9'd439},
      '{9'd007, 9'd014, 9'd028, 9'd056}, '{9'd263, 9'd015, 9'd029, 9'd057}, '{9'd135, 9'd270, 9'd030, 9'd058}, '{9'd391, 9'd271, 9'd031, 9'd059}, '{9'd071, 9'd142, 9'd284, 9'd060}, '{9'd327, 9'd143, 9'd285, 9'd061}, '{9'd199, 9'd398, 9'd286, 9'd062}, '{9'd455, 9'd399, 9'd287, 9'd063},
      '{9'd023, 9'd046, 9'd092, 9'd184}, '{9'd279, 9'd047, 9'd093, 9'd185}, '{9'd151, 9'd302, 9'd094, 9'd186}, '{9'd407, 9'd303, 9'd095, 9'd187}, '{9'd087, 9'd174, 9'd348, 9'd188}, '{9'd343, 9'd175, 9'd349, 9'd189}, '{9'd215, 9'd430, 9'd350, 9'd190}, '{9'd471, 9'd431, 9'd351, 9'd191},
      '{9'd039, 9'd078, 9'd156, 9'd312}, '{9'd295, 9'd079, 9'd157, 9'd313}, '{9'd167, 9'd334, 9'd158, 9'd314}, '{9'd423, 9'd335, 9'd159, 9'd315}, '{9'd103, 9'd206, 9'd412, 9'd316}, '{9'd359, 9'd207, 9'd413, 9'd317}, '{9'd231, 9'd462, 9'd414, 9'd318}, '{9'd487, 9'd463, 9'd415, 9'd319},
      '{9'd055, 9'd110, 9'd220, 9'd440}, '{9'd311, 9'd111, 9'd221, 9'd441}, '{9'd183, 9'd366, 9'd222, 9'd442}, '{9'd439, 9'd367, 9'd223, 9'd443}, '{9'd119, 9'd238, 9'd476, 9'd444}, '{9'd375, 9'd239, 9'd477, 9'd445}, '{9'd247, 9'd494, 9'd478, 9'd446}, '{9'd503, 9'd495, 9'd479, 9'd447},
      '{9'd008, 9'd016, 9'd032, 9'd064}, '{9'd264, 9'd017, 9'd033, 9'd065}, '{9'd136, 9'd272, 9'd034, 9'd066}, '{9'd392, 9'd273, 9'd035, 9'd067}, '{9'd072, 9'd144, 9'd288, 9'd068}, '{9'd328, 9'd145, 9'd289, 9'd069}, '{9'd200, 9'd400, 9'd290, 9'd070}, '{9'd456, 9'd401, 9'd291, 9'd071},
      '{9'd024, 9'd048, 9'd096, 9'd192}, '{9'd280, 9'd049, 9'd097, 9'd193}, '{9'd152, 9'd304, 9'd098, 9'd194}, '{9'd408, 9'd305, 9'd099, 9'd195}, '{9'd088, 9'd176, 9'd352, 9'd196}, '{9'd344, 9'd177, 9'd353, 9'd197}, '{9'd216, 9'd432, 9'd354, 9'd198}, '{9'd472, 9'd433, 9'd355, 9'd199},
      '{9'd040, 9'd080, 9'd160, 9'd320}, '{9'd296, 9'd081, 9'd161, 9'd321}, '{9'd168, 9'd336, 9'd162, 9'd322}, '{9'd424, 9'd337, 9'd163, 9'd323}, '{9'd104, 9'd208, 9'd416, 9'd324}, '{9'd360, 9'd209, 9'd417, 9'd325}, '{9'd232, 9'd464, 9'd418, 9'd326}, '{9'd488, 9'd465, 9'd419, 9'd327},
      '{9'd056, 9'd112, 9'd224, 9'd448}, '{9'd312, 9'd113, 9'd225, 9'd449}, '{9'd184, 9'd368, 9'd226, 9'd450}, '{9'd440, 9'd369, 9'd227, 9'd451}, '{9'd120, 9'd240, 9'd480, 9'd452}, '{9'd376, 9'd241, 9'd481, 9'd453}, '{9'd248, 9'd496, 9'd482, 9'd454}, '{9'd504, 9'd497, 9'd483, 9'd455},
      '{9'd009, 9'd018, 9'd036, 9'd072}, '{9'd265, 9'd019, 9'd037, 9'd073}, '{9'd137, 9'd274, 9'd038, 9'd074}, '{9'd393, 9'd275, 9'd039, 9'd075}, '{9'd073, 9'd146, 9'd292, 9'd076}, '{9'd329, 9'd147, 9'd293, 9'd077}, '{9'd201, 9'd402, 9'd294, 9'd078}, '{9'd457, 9'd403, 9'd295, 9'd079},
      '{9'd025, 9'd050, 9'd100, 9'd200}, '{9'd281, 9'd051, 9'd101, 9'd201}, '{9'd153, 9'd306, 9'd102, 9'd202}, '{9'd409, 9'd307, 9'd103, 9'd203}, '{9'd089, 9'd178, 9'd356, 9'd204}, '{9'd345, 9'd179, 9'd357, 9'd205}, '{9'd217, 9'd434, 9'd358, 9'd206}, '{9'd473, 9'd435, 9'd359, 9'd207},
      '{9'd041, 9'd082, 9'd164, 9'd328}, '{9'd297, 9'd083, 9'd165, 9'd329}, '{9'd169, 9'd338, 9'd166, 9'd330}, '{9'd425, 9'd339, 9'd167, 9'd331}, '{9'd105, 9'd210, 9'd420, 9'd332}, '{9'd361, 9'd211, 9'd421, 9'd333}, '{9'd233, 9'd466, 9'd422, 9'd334}, '{9'd489, 9'd467, 9'd423, 9'd335},
      '{9'd057, 9'd114, 9'd228, 9'd456}, '{9'd313, 9'd115, 9'd229, 9'd457}, '{9'd185, 9'd370, 9'd230, 9'd458}, '{9'd441, 9'd371, 9'd231, 9'd459}, '{9'd121, 9'd242, 9'd484, 9'd460}, '{9'd377, 9'd243, 9'd485, 9'd461}, '{9'd249, 9'd498, 9'd486, 9'd462}, '{9'd505, 9'd499, 9'd487, 9'd463},
      '{9'd010, 9'd020, 9'd040, 9'd080}, '{9'd266, 9'd021, 9'd041, 9'd081}, '{9'd138, 9'd276, 9'd042, 9'd082}, '{9'd394, 9'd277, 9'd043, 9'd083}, '{9'd074, 9'd148, 9'd296, 9'd084}, '{9'd330, 9'd149, 9'd297, 9'd085}, '{9'd202, 9'd404, 9'd298, 9'd086}, '{9'd458, 9'd405, 9'd299, 9'd087},
      '{9'd026, 9'd052, 9'd104, 9'd208}, '{9'd282, 9'd053, 9'd105, 9'd209}, '{9'd154, 9'd308, 9'd106, 9'd210}, '{9'd410, 9'd309, 9'd107, 9'd211}, '{9'd090, 9'd180, 9'd360, 9'd212}, '{9'd346, 9'd181, 9'd361, 9'd213}, '{9'd218, 9'd436, 9'd362, 9'd214}, '{9'd474, 9'd437, 9'd363, 9'd215},
      '{9'd042, 9'd084, 9'd168, 9'd336}, '{9'd298, 9'd085, 9'd169, 9'd337}, '{9'd170, 9'd340, 9'd170, 9'd338}, '{9'd426, 9'd341, 9'd171, 9'd339}, '{9'd106, 9'd212, 9'd424, 9'd340}, '{9'd362, 9'd213, 9'd425, 9'd341}, '{9'd234, 9'd468, 9'd426, 9'd342}, '{9'd490, 9'd469, 9'd427, 9'd343},
      '{9'd058, 9'd116, 9'd232, 9'd464}, '{9'd314, 9'd117, 9'd233, 9'd465}, '{9'd186, 9'd372, 9'd234, 9'd466}, '{9'd442, 9'd373, 9'd235, 9'd467}, '{9'd122, 9'd244, 9'd488, 9'd468}, '{9'd378, 9'd245, 9'd489, 9'd469}, '{9'd250, 9'd500, 9'd490, 9'd470}, '{9'd506, 9'd501, 9'd491, 9'd471},
      '{9'd011, 9'd022, 9'd044, 9'd088}, '{9'd267, 9'd023, 9'd045, 9'd089}, '{9'd139, 9'd278, 9'd046, 9'd090}, '{9'd395, 9'd279, 9'd047, 9'd091}, '{9'd075, 9'd150, 9'd300, 9'd092}, '{9'd331, 9'd151, 9'd301, 9'd093}, '{9'd203, 9'd406, 9'd302, 9'd094}, '{9'd459, 9'd407, 9'd303, 9'd095},
      '{9'd027, 9'd054, 9'd108, 9'd216}, '{9'd283, 9'd055, 9'd109, 9'd217}, '{9'd155, 9'd310, 9'd110, 9'd218}, '{9'd411, 9'd311, 9'd111, 9'd219}, '{9'd091, 9'd182, 9'd364, 9'd220}, '{9'd347, 9'd183, 9'd365, 9'd221}, '{9'd219, 9'd438, 9'd366, 9'd222}, '{9'd475, 9'd439, 9'd367, 9'd223},
      '{9'd043, 9'd086, 9'd172, 9'd344}, '{9'd299, 9'd087, 9'd173, 9'd345}, '{9'd171, 9'd342, 9'd174, 9'd346}, '{9'd427, 9'd343, 9'd175, 9'd347}, '{9'd107, 9'd214, 9'd428, 9'd348}, '{9'd363, 9'd215, 9'd429, 9'd349}, '{9'd235, 9'd470, 9'd430, 9'd350}, '{9'd491, 9'd471, 9'd431, 9'd351},
      '{9'd059, 9'd118, 9'd236, 9'd472}, '{9'd315, 9'd119, 9'd237, 9'd473}, '{9'd187, 9'd374, 9'd238, 9'd474}, '{9'd443, 9'd375, 9'd239, 9'd475}, '{9'd123, 9'd246, 9'd492, 9'd476}, '{9'd379, 9'd247, 9'd493, 9'd477}, '{9'd251, 9'd502, 9'd494, 9'd478}, '{9'd507, 9'd503, 9'd495, 9'd479},
      '{9'd012, 9'd024, 9'd048, 9'd096}, '{9'd268, 9'd025, 9'd049, 9'd097}, '{9'd140, 9'd280, 9'd050, 9'd098}, '{9'd396, 9'd281, 9'd051, 9'd099}, '{9'd076, 9'd152, 9'd304, 9'd100}, '{9'd332, 9'd153, 9'd305, 9'd101}, '{9'd204, 9'd408, 9'd306, 9'd102}, '{9'd460, 9'd409, 9'd307, 9'd103},
      '{9'd028, 9'd056, 9'd112, 9'd224}, '{9'd284, 9'd057, 9'd113, 9'd225}, '{9'd156, 9'd312, 9'd114, 9'd226}, '{9'd412, 9'd313, 9'd115, 9'd227}, '{9'd092, 9'd184, 9'd368, 9'd228}, '{9'd348, 9'd185, 9'd369, 9'd229}, '{9'd220, 9'd440, 9'd370, 9'd230}, '{9'd476, 9'd441, 9'd371, 9'd231},
      '{9'd044, 9'd088, 9'd176, 9'd352}, '{9'd300, 9'd089, 9'd177, 9'd353}, '{9'd172, 9'd344, 9'd178, 9'd354}, '{9'd428, 9'd345, 9'd179, 9'd355}, '{9'd108, 9'd216, 9'd432, 9'd356}, '{9'd364, 9'd217, 9'd433, 9'd357}, '{9'd236, 9'd472, 9'd434, 9'd358}, '{9'd492, 9'd473, 9'd435, 9'd359},
      '{9'd060, 9'd120, 9'd240, 9'd480}, '{9'd316, 9'd121, 9'd241, 9'd481}, '{9'd188, 9'd376, 9'd242, 9'd482}, '{9'd444, 9'd377, 9'd243, 9'd483}, '{9'd124, 9'd248, 9'd496, 9'd484}, '{9'd380, 9'd249, 9'd497, 9'd485}, '{9'd252, 9'd504, 9'd498, 9'd486}, '{9'd508, 9'd505, 9'd499, 9'd487},
      '{9'd013, 9'd026, 9'd052, 9'd104}, '{9'd269, 9'd027, 9'd053, 9'd105}, '{9'd141, 9'd282, 9'd054, 9'd106}, '{9'd397, 9'd283, 9'd055, 9'd107}, '{9'd077, 9'd154, 9'd308, 9'd108}, '{9'd333, 9'd155, 9'd309, 9'd109}, '{9'd205, 9'd410, 9'd310, 9'd110}, '{9'd461, 9'd411, 9'd311, 9'd111},
      '{9'd029, 9'd058, 9'd116, 9'd232}, '{9'd285, 9'd059, 9'd117, 9'd233}, '{9'd157, 9'd314, 9'd118, 9'd234}, '{9'd413, 9'd315, 9'd119, 9'd235}, '{9'd093, 9'd186, 9'd372, 9'd236}, '{9'd349, 9'd187, 9'd373, 9'd237}, '{9'd221, 9'd442, 9'd374, 9'd238}, '{9'd477, 9'd443, 9'd375, 9'd239},
      '{9'd045, 9'd090, 9'd180, 9'd360}, '{9'd301, 9'd091, 9'd181, 9'd361}, '{9'd173, 9'd346, 9'd182, 9'd362}, '{9'd429, 9'd347, 9'd183, 9'd363}, '{9'd109, 9'd218, 9'd436, 9'd364}, '{9'd365, 9'd219, 9'd437, 9'd365}, '{9'd237, 9'd474, 9'd438, 9'd366}, '{9'd493, 9'd475, 9'd439, 9'd367},
      '{9'd061, 9'd122, 9'd244, 9'd488}, '{9'd317, 9'd123, 9'd245, 9'd489}, '{9'd189, 9'd378, 9'd246, 9'd490}, '{9'd445, 9'd379, 9'd247, 9'd491}, '{9'd125, 9'd250, 9'd500, 9'd492}, '{9'd381, 9'd251, 9'd501, 9'd493}, '{9'd253, 9'd506, 9'd502, 9'd494}, '{9'd509, 9'd507, 9'd503, 9'd495},
      '{9'd014, 9'd028, 9'd056, 9'd112}, '{9'd270, 9'd029, 9'd057, 9'd113}, '{9'd142, 9'd284, 9'd058, 9'd114}, '{9'd398, 9'd285, 9'd059, 9'd115}, '{9'd078, 9'd156, 9'd312, 9'd116}, '{9'd334, 9'd157, 9'd313, 9'd117}, '{9'd206, 9'd412, 9'd314, 9'd118}, '{9'd462, 9'd413, 9'd315, 9'd119},
      '{9'd030, 9'd060, 9'd120, 9'd240}, '{9'd286, 9'd061, 9'd121, 9'd241}, '{9'd158, 9'd316, 9'd122, 9'd242}, '{9'd414, 9'd317, 9'd123, 9'd243}, '{9'd094, 9'd188, 9'd376, 9'd244}, '{9'd350, 9'd189, 9'd377, 9'd245}, '{9'd222, 9'd444, 9'd378, 9'd246}, '{9'd478, 9'd445, 9'd379, 9'd247},
      '{9'd046, 9'd092, 9'd184, 9'd368}, '{9'd302, 9'd093, 9'd185, 9'd369}, '{9'd174, 9'd348, 9'd186, 9'd370}, '{9'd430, 9'd349, 9'd187, 9'd371}, '{9'd110, 9'd220, 9'd440, 9'd372}, '{9'd366, 9'd221, 9'd441, 9'd373}, '{9'd238, 9'd476, 9'd442, 9'd374}, '{9'd494, 9'd477, 9'd443, 9'd375},
      '{9'd062, 9'd124, 9'd248, 9'd496}, '{9'd318, 9'd125, 9'd249, 9'd497}, '{9'd190, 9'd380, 9'd250, 9'd498}, '{9'd446, 9'd381, 9'd251, 9'd499}, '{9'd126, 9'd252, 9'd504, 9'd500}, '{9'd382, 9'd253, 9'd505, 9'd501}, '{9'd254, 9'd508, 9'd506, 9'd502}, '{9'd510, 9'd509, 9'd507, 9'd503},
      '{9'd015, 9'd030, 9'd060, 9'd120}, '{9'd271, 9'd031, 9'd061, 9'd121}, '{9'd143, 9'd286, 9'd062, 9'd122}, '{9'd399, 9'd287, 9'd063, 9'd123}, '{9'd079, 9'd158, 9'd316, 9'd124}, '{9'd335, 9'd159, 9'd317, 9'd125}, '{9'd207, 9'd414, 9'd318, 9'd126}, '{9'd463, 9'd415, 9'd319, 9'd127},
      '{9'd031, 9'd062, 9'd124, 9'd248}, '{9'd287, 9'd063, 9'd125, 9'd249}, '{9'd159, 9'd318, 9'd126, 9'd250}, '{9'd415, 9'd319, 9'd127, 9'd251}, '{9'd095, 9'd190, 9'd380, 9'd252}, '{9'd351, 9'd191, 9'd381, 9'd253}, '{9'd223, 9'd446, 9'd382, 9'd254}, '{9'd479, 9'd447, 9'd383, 9'd255},
      '{9'd047, 9'd094, 9'd188, 9'd376}, '{9'd303, 9'd095, 9'd189, 9'd377}, '{9'd175, 9'd350, 9'd190, 9'd378}, '{9'd431, 9'd351, 9'd191, 9'd379}, '{9'd111, 9'd222, 9'd444, 9'd380}, '{9'd367, 9'd223, 9'd445, 9'd381}, '{9'd239, 9'd478, 9'd446, 9'd382}, '{9'd495, 9'd479, 9'd447, 9'd383},
      '{9'd063, 9'd126, 9'd252, 9'd504}, '{9'd319, 9'd127, 9'd253, 9'd505}, '{9'd191, 9'd382, 9'd254, 9'd506}, '{9'd447, 9'd383, 9'd255, 9'd507}, '{9'd127, 9'd254, 9'd508, 9'd508}, '{9'd383, 9'd255, 9'd509, 9'd509}, '{9'd255, 9'd510, 9'd510, 9'd510}, '{9'd511, 9'd511, 9'd511, 9'd511}
    };

    unique case (NrLanes)
      1 : return lut_1lane [shfNbIdx][ew];
      2 : return lut_2lane [shfNbIdx][ew];
      4 : return lut_4lane [shfNbIdx][ew];
      8 : return lut_8lane [shfNbIdx][ew];
      16: return lut_16lane[shfNbIdx][ew];
      default: return 0;
	  endcase
  endfunction

  function automatic logic [{$clog2(riva_pkg::DLEN*riva_pkg::MaxNrLanes/4)}-1:0] query_seq_idx_2d_cln(input int NrLanes, input int shfNbIdx, input riscv_mv_pkg::vew_e ew);
    automatic logic [5-1:0] lut_1lane [0:31][0:3] = '{
      '{5'd000, 5'd000, 5'd000, 5'd000}, '{5'd016, 5'd001, 5'd001, 5'd001}, '{5'd008, 5'd016, 5'd002, 5'd002}, '{5'd024, 5'd017, 5'd003, 5'd003}, '{5'd004, 5'd008, 5'd016, 5'd004}, '{5'd020, 5'd009, 5'd017, 5'd005}, '{5'd012, 5'd024, 5'd018, 5'd006}, '{5'd028, 5'd025, 5'd019, 5'd007},
      '{5'd001, 5'd002, 5'd004, 5'd008}, '{5'd017, 5'd003, 5'd005, 5'd009}, '{5'd009, 5'd018, 5'd006, 5'd010}, '{5'd025, 5'd019, 5'd007, 5'd011}, '{5'd005, 5'd010, 5'd020, 5'd012}, '{5'd021, 5'd011, 5'd021, 5'd013}, '{5'd013, 5'd026, 5'd022, 5'd014}, '{5'd029, 5'd027, 5'd023, 5'd015},
      '{5'd002, 5'd004, 5'd008, 5'd016}, '{5'd018, 5'd005, 5'd009, 5'd017}, '{5'd010, 5'd020, 5'd010, 5'd018}, '{5'd026, 5'd021, 5'd011, 5'd019}, '{5'd006, 5'd012, 5'd024, 5'd020}, '{5'd022, 5'd013, 5'd025, 5'd021}, '{5'd014, 5'd028, 5'd026, 5'd022}, '{5'd030, 5'd029, 5'd027, 5'd023},
      '{5'd003, 5'd006, 5'd012, 5'd024}, '{5'd019, 5'd007, 5'd013, 5'd025}, '{5'd011, 5'd022, 5'd014, 5'd026}, '{5'd027, 5'd023, 5'd015, 5'd027}, '{5'd007, 5'd014, 5'd028, 5'd028}, '{5'd023, 5'd015, 5'd029, 5'd029}, '{5'd015, 5'd030, 5'd030, 5'd030}, '{5'd031, 5'd031, 5'd031, 5'd031}
    };
    automatic logic [6-1:0] lut_2lane [0:63][0:3] = '{
      '{6'd000, 6'd000, 6'd000, 6'd000}, '{6'd016, 6'd001, 6'd001, 6'd001}, '{6'd008, 6'd016, 6'd002, 6'd002}, '{6'd024, 6'd017, 6'd003, 6'd003}, '{6'd004, 6'd008, 6'd016, 6'd004}, '{6'd020, 6'd009, 6'd017, 6'd005}, '{6'd012, 6'd024, 6'd018, 6'd006}, '{6'd028, 6'd025, 6'd019, 6'd007},
      '{6'd001, 6'd002, 6'd004, 6'd008}, '{6'd017, 6'd003, 6'd005, 6'd009}, '{6'd009, 6'd018, 6'd006, 6'd010}, '{6'd025, 6'd019, 6'd007, 6'd011}, '{6'd005, 6'd010, 6'd020, 6'd012}, '{6'd021, 6'd011, 6'd021, 6'd013}, '{6'd013, 6'd026, 6'd022, 6'd014}, '{6'd029, 6'd027, 6'd023, 6'd015},
      '{6'd002, 6'd004, 6'd008, 6'd016}, '{6'd018, 6'd005, 6'd009, 6'd017}, '{6'd010, 6'd020, 6'd010, 6'd018}, '{6'd026, 6'd021, 6'd011, 6'd019}, '{6'd006, 6'd012, 6'd024, 6'd020}, '{6'd022, 6'd013, 6'd025, 6'd021}, '{6'd014, 6'd028, 6'd026, 6'd022}, '{6'd030, 6'd029, 6'd027, 6'd023},
      '{6'd003, 6'd006, 6'd012, 6'd024}, '{6'd019, 6'd007, 6'd013, 6'd025}, '{6'd011, 6'd022, 6'd014, 6'd026}, '{6'd027, 6'd023, 6'd015, 6'd027}, '{6'd007, 6'd014, 6'd028, 6'd028}, '{6'd023, 6'd015, 6'd029, 6'd029}, '{6'd015, 6'd030, 6'd030, 6'd030}, '{6'd031, 6'd031, 6'd031, 6'd031},
      '{6'd032, 6'd032, 6'd032, 6'd032}, '{6'd048, 6'd033, 6'd033, 6'd033}, '{6'd040, 6'd048, 6'd034, 6'd034}, '{6'd056, 6'd049, 6'd035, 6'd035}, '{6'd036, 6'd040, 6'd048, 6'd036}, '{6'd052, 6'd041, 6'd049, 6'd037}, '{6'd044, 6'd056, 6'd050, 6'd038}, '{6'd060, 6'd057, 6'd051, 6'd039},
      '{6'd033, 6'd034, 6'd036, 6'd040}, '{6'd049, 6'd035, 6'd037, 6'd041}, '{6'd041, 6'd050, 6'd038, 6'd042}, '{6'd057, 6'd051, 6'd039, 6'd043}, '{6'd037, 6'd042, 6'd052, 6'd044}, '{6'd053, 6'd043, 6'd053, 6'd045}, '{6'd045, 6'd058, 6'd054, 6'd046}, '{6'd061, 6'd059, 6'd055, 6'd047},
      '{6'd034, 6'd036, 6'd040, 6'd048}, '{6'd050, 6'd037, 6'd041, 6'd049}, '{6'd042, 6'd052, 6'd042, 6'd050}, '{6'd058, 6'd053, 6'd043, 6'd051}, '{6'd038, 6'd044, 6'd056, 6'd052}, '{6'd054, 6'd045, 6'd057, 6'd053}, '{6'd046, 6'd060, 6'd058, 6'd054}, '{6'd062, 6'd061, 6'd059, 6'd055},
      '{6'd035, 6'd038, 6'd044, 6'd056}, '{6'd051, 6'd039, 6'd045, 6'd057}, '{6'd043, 6'd054, 6'd046, 6'd058}, '{6'd059, 6'd055, 6'd047, 6'd059}, '{6'd039, 6'd046, 6'd060, 6'd060}, '{6'd055, 6'd047, 6'd061, 6'd061}, '{6'd047, 6'd062, 6'd062, 6'd062}, '{6'd063, 6'd063, 6'd063, 6'd063}
    };
    automatic logic [7-1:0] lut_4lane [0:127][0:3] = '{
      '{7'd000, 7'd000, 7'd000, 7'd000}, '{7'd016, 7'd001, 7'd001, 7'd001}, '{7'd008, 7'd016, 7'd002, 7'd002}, '{7'd024, 7'd017, 7'd003, 7'd003}, '{7'd004, 7'd008, 7'd016, 7'd004}, '{7'd020, 7'd009, 7'd017, 7'd005}, '{7'd012, 7'd024, 7'd018, 7'd006}, '{7'd028, 7'd025, 7'd019, 7'd007},
      '{7'd001, 7'd002, 7'd004, 7'd008}, '{7'd017, 7'd003, 7'd005, 7'd009}, '{7'd009, 7'd018, 7'd006, 7'd010}, '{7'd025, 7'd019, 7'd007, 7'd011}, '{7'd005, 7'd010, 7'd020, 7'd012}, '{7'd021, 7'd011, 7'd021, 7'd013}, '{7'd013, 7'd026, 7'd022, 7'd014}, '{7'd029, 7'd027, 7'd023, 7'd015},
      '{7'd002, 7'd004, 7'd008, 7'd016}, '{7'd018, 7'd005, 7'd009, 7'd017}, '{7'd010, 7'd020, 7'd010, 7'd018}, '{7'd026, 7'd021, 7'd011, 7'd019}, '{7'd006, 7'd012, 7'd024, 7'd020}, '{7'd022, 7'd013, 7'd025, 7'd021}, '{7'd014, 7'd028, 7'd026, 7'd022}, '{7'd030, 7'd029, 7'd027, 7'd023},
      '{7'd003, 7'd006, 7'd012, 7'd024}, '{7'd019, 7'd007, 7'd013, 7'd025}, '{7'd011, 7'd022, 7'd014, 7'd026}, '{7'd027, 7'd023, 7'd015, 7'd027}, '{7'd007, 7'd014, 7'd028, 7'd028}, '{7'd023, 7'd015, 7'd029, 7'd029}, '{7'd015, 7'd030, 7'd030, 7'd030}, '{7'd031, 7'd031, 7'd031, 7'd031},
      '{7'd032, 7'd032, 7'd032, 7'd032}, '{7'd048, 7'd033, 7'd033, 7'd033}, '{7'd040, 7'd048, 7'd034, 7'd034}, '{7'd056, 7'd049, 7'd035, 7'd035}, '{7'd036, 7'd040, 7'd048, 7'd036}, '{7'd052, 7'd041, 7'd049, 7'd037}, '{7'd044, 7'd056, 7'd050, 7'd038}, '{7'd060, 7'd057, 7'd051, 7'd039},
      '{7'd033, 7'd034, 7'd036, 7'd040}, '{7'd049, 7'd035, 7'd037, 7'd041}, '{7'd041, 7'd050, 7'd038, 7'd042}, '{7'd057, 7'd051, 7'd039, 7'd043}, '{7'd037, 7'd042, 7'd052, 7'd044}, '{7'd053, 7'd043, 7'd053, 7'd045}, '{7'd045, 7'd058, 7'd054, 7'd046}, '{7'd061, 7'd059, 7'd055, 7'd047},
      '{7'd034, 7'd036, 7'd040, 7'd048}, '{7'd050, 7'd037, 7'd041, 7'd049}, '{7'd042, 7'd052, 7'd042, 7'd050}, '{7'd058, 7'd053, 7'd043, 7'd051}, '{7'd038, 7'd044, 7'd056, 7'd052}, '{7'd054, 7'd045, 7'd057, 7'd053}, '{7'd046, 7'd060, 7'd058, 7'd054}, '{7'd062, 7'd061, 7'd059, 7'd055},
      '{7'd035, 7'd038, 7'd044, 7'd056}, '{7'd051, 7'd039, 7'd045, 7'd057}, '{7'd043, 7'd054, 7'd046, 7'd058}, '{7'd059, 7'd055, 7'd047, 7'd059}, '{7'd039, 7'd046, 7'd060, 7'd060}, '{7'd055, 7'd047, 7'd061, 7'd061}, '{7'd047, 7'd062, 7'd062, 7'd062}, '{7'd063, 7'd063, 7'd063, 7'd063},
      '{7'd064, 7'd064, 7'd064, 7'd064}, '{7'd080, 7'd065, 7'd065, 7'd065}, '{7'd072, 7'd080, 7'd066, 7'd066}, '{7'd088, 7'd081, 7'd067, 7'd067}, '{7'd068, 7'd072, 7'd080, 7'd068}, '{7'd084, 7'd073, 7'd081, 7'd069}, '{7'd076, 7'd088, 7'd082, 7'd070}, '{7'd092, 7'd089, 7'd083, 7'd071},
      '{7'd065, 7'd066, 7'd068, 7'd072}, '{7'd081, 7'd067, 7'd069, 7'd073}, '{7'd073, 7'd082, 7'd070, 7'd074}, '{7'd089, 7'd083, 7'd071, 7'd075}, '{7'd069, 7'd074, 7'd084, 7'd076}, '{7'd085, 7'd075, 7'd085, 7'd077}, '{7'd077, 7'd090, 7'd086, 7'd078}, '{7'd093, 7'd091, 7'd087, 7'd079},
      '{7'd066, 7'd068, 7'd072, 7'd080}, '{7'd082, 7'd069, 7'd073, 7'd081}, '{7'd074, 7'd084, 7'd074, 7'd082}, '{7'd090, 7'd085, 7'd075, 7'd083}, '{7'd070, 7'd076, 7'd088, 7'd084}, '{7'd086, 7'd077, 7'd089, 7'd085}, '{7'd078, 7'd092, 7'd090, 7'd086}, '{7'd094, 7'd093, 7'd091, 7'd087},
      '{7'd067, 7'd070, 7'd076, 7'd088}, '{7'd083, 7'd071, 7'd077, 7'd089}, '{7'd075, 7'd086, 7'd078, 7'd090}, '{7'd091, 7'd087, 7'd079, 7'd091}, '{7'd071, 7'd078, 7'd092, 7'd092}, '{7'd087, 7'd079, 7'd093, 7'd093}, '{7'd079, 7'd094, 7'd094, 7'd094}, '{7'd095, 7'd095, 7'd095, 7'd095},
      '{7'd096, 7'd096, 7'd096, 7'd096}, '{7'd112, 7'd097, 7'd097, 7'd097}, '{7'd104, 7'd112, 7'd098, 7'd098}, '{7'd120, 7'd113, 7'd099, 7'd099}, '{7'd100, 7'd104, 7'd112, 7'd100}, '{7'd116, 7'd105, 7'd113, 7'd101}, '{7'd108, 7'd120, 7'd114, 7'd102}, '{7'd124, 7'd121, 7'd115, 7'd103},
      '{7'd097, 7'd098, 7'd100, 7'd104}, '{7'd113, 7'd099, 7'd101, 7'd105}, '{7'd105, 7'd114, 7'd102, 7'd106}, '{7'd121, 7'd115, 7'd103, 7'd107}, '{7'd101, 7'd106, 7'd116, 7'd108}, '{7'd117, 7'd107, 7'd117, 7'd109}, '{7'd109, 7'd122, 7'd118, 7'd110}, '{7'd125, 7'd123, 7'd119, 7'd111},
      '{7'd098, 7'd100, 7'd104, 7'd112}, '{7'd114, 7'd101, 7'd105, 7'd113}, '{7'd106, 7'd116, 7'd106, 7'd114}, '{7'd122, 7'd117, 7'd107, 7'd115}, '{7'd102, 7'd108, 7'd120, 7'd116}, '{7'd118, 7'd109, 7'd121, 7'd117}, '{7'd110, 7'd124, 7'd122, 7'd118}, '{7'd126, 7'd125, 7'd123, 7'd119},
      '{7'd099, 7'd102, 7'd108, 7'd120}, '{7'd115, 7'd103, 7'd109, 7'd121}, '{7'd107, 7'd118, 7'd110, 7'd122}, '{7'd123, 7'd119, 7'd111, 7'd123}, '{7'd103, 7'd110, 7'd124, 7'd124}, '{7'd119, 7'd111, 7'd125, 7'd125}, '{7'd111, 7'd126, 7'd126, 7'd126}, '{7'd127, 7'd127, 7'd127, 7'd127}
    };
    automatic logic [8-1:0] lut_8lane [0:255][0:3] = '{
      '{8'd000, 8'd000, 8'd000, 8'd000}, '{8'd016, 8'd001, 8'd001, 8'd001}, '{8'd008, 8'd016, 8'd002, 8'd002}, '{8'd024, 8'd017, 8'd003, 8'd003}, '{8'd004, 8'd008, 8'd016, 8'd004}, '{8'd020, 8'd009, 8'd017, 8'd005}, '{8'd012, 8'd024, 8'd018, 8'd006}, '{8'd028, 8'd025, 8'd019, 8'd007},
      '{8'd001, 8'd002, 8'd004, 8'd008}, '{8'd017, 8'd003, 8'd005, 8'd009}, '{8'd009, 8'd018, 8'd006, 8'd010}, '{8'd025, 8'd019, 8'd007, 8'd011}, '{8'd005, 8'd010, 8'd020, 8'd012}, '{8'd021, 8'd011, 8'd021, 8'd013}, '{8'd013, 8'd026, 8'd022, 8'd014}, '{8'd029, 8'd027, 8'd023, 8'd015},
      '{8'd002, 8'd004, 8'd008, 8'd016}, '{8'd018, 8'd005, 8'd009, 8'd017}, '{8'd010, 8'd020, 8'd010, 8'd018}, '{8'd026, 8'd021, 8'd011, 8'd019}, '{8'd006, 8'd012, 8'd024, 8'd020}, '{8'd022, 8'd013, 8'd025, 8'd021}, '{8'd014, 8'd028, 8'd026, 8'd022}, '{8'd030, 8'd029, 8'd027, 8'd023},
      '{8'd003, 8'd006, 8'd012, 8'd024}, '{8'd019, 8'd007, 8'd013, 8'd025}, '{8'd011, 8'd022, 8'd014, 8'd026}, '{8'd027, 8'd023, 8'd015, 8'd027}, '{8'd007, 8'd014, 8'd028, 8'd028}, '{8'd023, 8'd015, 8'd029, 8'd029}, '{8'd015, 8'd030, 8'd030, 8'd030}, '{8'd031, 8'd031, 8'd031, 8'd031},
      '{8'd032, 8'd032, 8'd032, 8'd032}, '{8'd048, 8'd033, 8'd033, 8'd033}, '{8'd040, 8'd048, 8'd034, 8'd034}, '{8'd056, 8'd049, 8'd035, 8'd035}, '{8'd036, 8'd040, 8'd048, 8'd036}, '{8'd052, 8'd041, 8'd049, 8'd037}, '{8'd044, 8'd056, 8'd050, 8'd038}, '{8'd060, 8'd057, 8'd051, 8'd039},
      '{8'd033, 8'd034, 8'd036, 8'd040}, '{8'd049, 8'd035, 8'd037, 8'd041}, '{8'd041, 8'd050, 8'd038, 8'd042}, '{8'd057, 8'd051, 8'd039, 8'd043}, '{8'd037, 8'd042, 8'd052, 8'd044}, '{8'd053, 8'd043, 8'd053, 8'd045}, '{8'd045, 8'd058, 8'd054, 8'd046}, '{8'd061, 8'd059, 8'd055, 8'd047},
      '{8'd034, 8'd036, 8'd040, 8'd048}, '{8'd050, 8'd037, 8'd041, 8'd049}, '{8'd042, 8'd052, 8'd042, 8'd050}, '{8'd058, 8'd053, 8'd043, 8'd051}, '{8'd038, 8'd044, 8'd056, 8'd052}, '{8'd054, 8'd045, 8'd057, 8'd053}, '{8'd046, 8'd060, 8'd058, 8'd054}, '{8'd062, 8'd061, 8'd059, 8'd055},
      '{8'd035, 8'd038, 8'd044, 8'd056}, '{8'd051, 8'd039, 8'd045, 8'd057}, '{8'd043, 8'd054, 8'd046, 8'd058}, '{8'd059, 8'd055, 8'd047, 8'd059}, '{8'd039, 8'd046, 8'd060, 8'd060}, '{8'd055, 8'd047, 8'd061, 8'd061}, '{8'd047, 8'd062, 8'd062, 8'd062}, '{8'd063, 8'd063, 8'd063, 8'd063},
      '{8'd064, 8'd064, 8'd064, 8'd064}, '{8'd080, 8'd065, 8'd065, 8'd065}, '{8'd072, 8'd080, 8'd066, 8'd066}, '{8'd088, 8'd081, 8'd067, 8'd067}, '{8'd068, 8'd072, 8'd080, 8'd068}, '{8'd084, 8'd073, 8'd081, 8'd069}, '{8'd076, 8'd088, 8'd082, 8'd070}, '{8'd092, 8'd089, 8'd083, 8'd071},
      '{8'd065, 8'd066, 8'd068, 8'd072}, '{8'd081, 8'd067, 8'd069, 8'd073}, '{8'd073, 8'd082, 8'd070, 8'd074}, '{8'd089, 8'd083, 8'd071, 8'd075}, '{8'd069, 8'd074, 8'd084, 8'd076}, '{8'd085, 8'd075, 8'd085, 8'd077}, '{8'd077, 8'd090, 8'd086, 8'd078}, '{8'd093, 8'd091, 8'd087, 8'd079},
      '{8'd066, 8'd068, 8'd072, 8'd080}, '{8'd082, 8'd069, 8'd073, 8'd081}, '{8'd074, 8'd084, 8'd074, 8'd082}, '{8'd090, 8'd085, 8'd075, 8'd083}, '{8'd070, 8'd076, 8'd088, 8'd084}, '{8'd086, 8'd077, 8'd089, 8'd085}, '{8'd078, 8'd092, 8'd090, 8'd086}, '{8'd094, 8'd093, 8'd091, 8'd087},
      '{8'd067, 8'd070, 8'd076, 8'd088}, '{8'd083, 8'd071, 8'd077, 8'd089}, '{8'd075, 8'd086, 8'd078, 8'd090}, '{8'd091, 8'd087, 8'd079, 8'd091}, '{8'd071, 8'd078, 8'd092, 8'd092}, '{8'd087, 8'd079, 8'd093, 8'd093}, '{8'd079, 8'd094, 8'd094, 8'd094}, '{8'd095, 8'd095, 8'd095, 8'd095},
      '{8'd096, 8'd096, 8'd096, 8'd096}, '{8'd112, 8'd097, 8'd097, 8'd097}, '{8'd104, 8'd112, 8'd098, 8'd098}, '{8'd120, 8'd113, 8'd099, 8'd099}, '{8'd100, 8'd104, 8'd112, 8'd100}, '{8'd116, 8'd105, 8'd113, 8'd101}, '{8'd108, 8'd120, 8'd114, 8'd102}, '{8'd124, 8'd121, 8'd115, 8'd103},
      '{8'd097, 8'd098, 8'd100, 8'd104}, '{8'd113, 8'd099, 8'd101, 8'd105}, '{8'd105, 8'd114, 8'd102, 8'd106}, '{8'd121, 8'd115, 8'd103, 8'd107}, '{8'd101, 8'd106, 8'd116, 8'd108}, '{8'd117, 8'd107, 8'd117, 8'd109}, '{8'd109, 8'd122, 8'd118, 8'd110}, '{8'd125, 8'd123, 8'd119, 8'd111},
      '{8'd098, 8'd100, 8'd104, 8'd112}, '{8'd114, 8'd101, 8'd105, 8'd113}, '{8'd106, 8'd116, 8'd106, 8'd114}, '{8'd122, 8'd117, 8'd107, 8'd115}, '{8'd102, 8'd108, 8'd120, 8'd116}, '{8'd118, 8'd109, 8'd121, 8'd117}, '{8'd110, 8'd124, 8'd122, 8'd118}, '{8'd126, 8'd125, 8'd123, 8'd119},
      '{8'd099, 8'd102, 8'd108, 8'd120}, '{8'd115, 8'd103, 8'd109, 8'd121}, '{8'd107, 8'd118, 8'd110, 8'd122}, '{8'd123, 8'd119, 8'd111, 8'd123}, '{8'd103, 8'd110, 8'd124, 8'd124}, '{8'd119, 8'd111, 8'd125, 8'd125}, '{8'd111, 8'd126, 8'd126, 8'd126}, '{8'd127, 8'd127, 8'd127, 8'd127},
      '{8'd128, 8'd128, 8'd128, 8'd128}, '{8'd144, 8'd129, 8'd129, 8'd129}, '{8'd136, 8'd144, 8'd130, 8'd130}, '{8'd152, 8'd145, 8'd131, 8'd131}, '{8'd132, 8'd136, 8'd144, 8'd132}, '{8'd148, 8'd137, 8'd145, 8'd133}, '{8'd140, 8'd152, 8'd146, 8'd134}, '{8'd156, 8'd153, 8'd147, 8'd135},
      '{8'd129, 8'd130, 8'd132, 8'd136}, '{8'd145, 8'd131, 8'd133, 8'd137}, '{8'd137, 8'd146, 8'd134, 8'd138}, '{8'd153, 8'd147, 8'd135, 8'd139}, '{8'd133, 8'd138, 8'd148, 8'd140}, '{8'd149, 8'd139, 8'd149, 8'd141}, '{8'd141, 8'd154, 8'd150, 8'd142}, '{8'd157, 8'd155, 8'd151, 8'd143},
      '{8'd130, 8'd132, 8'd136, 8'd144}, '{8'd146, 8'd133, 8'd137, 8'd145}, '{8'd138, 8'd148, 8'd138, 8'd146}, '{8'd154, 8'd149, 8'd139, 8'd147}, '{8'd134, 8'd140, 8'd152, 8'd148}, '{8'd150, 8'd141, 8'd153, 8'd149}, '{8'd142, 8'd156, 8'd154, 8'd150}, '{8'd158, 8'd157, 8'd155, 8'd151},
      '{8'd131, 8'd134, 8'd140, 8'd152}, '{8'd147, 8'd135, 8'd141, 8'd153}, '{8'd139, 8'd150, 8'd142, 8'd154}, '{8'd155, 8'd151, 8'd143, 8'd155}, '{8'd135, 8'd142, 8'd156, 8'd156}, '{8'd151, 8'd143, 8'd157, 8'd157}, '{8'd143, 8'd158, 8'd158, 8'd158}, '{8'd159, 8'd159, 8'd159, 8'd159},
      '{8'd160, 8'd160, 8'd160, 8'd160}, '{8'd176, 8'd161, 8'd161, 8'd161}, '{8'd168, 8'd176, 8'd162, 8'd162}, '{8'd184, 8'd177, 8'd163, 8'd163}, '{8'd164, 8'd168, 8'd176, 8'd164}, '{8'd180, 8'd169, 8'd177, 8'd165}, '{8'd172, 8'd184, 8'd178, 8'd166}, '{8'd188, 8'd185, 8'd179, 8'd167},
      '{8'd161, 8'd162, 8'd164, 8'd168}, '{8'd177, 8'd163, 8'd165, 8'd169}, '{8'd169, 8'd178, 8'd166, 8'd170}, '{8'd185, 8'd179, 8'd167, 8'd171}, '{8'd165, 8'd170, 8'd180, 8'd172}, '{8'd181, 8'd171, 8'd181, 8'd173}, '{8'd173, 8'd186, 8'd182, 8'd174}, '{8'd189, 8'd187, 8'd183, 8'd175},
      '{8'd162, 8'd164, 8'd168, 8'd176}, '{8'd178, 8'd165, 8'd169, 8'd177}, '{8'd170, 8'd180, 8'd170, 8'd178}, '{8'd186, 8'd181, 8'd171, 8'd179}, '{8'd166, 8'd172, 8'd184, 8'd180}, '{8'd182, 8'd173, 8'd185, 8'd181}, '{8'd174, 8'd188, 8'd186, 8'd182}, '{8'd190, 8'd189, 8'd187, 8'd183},
      '{8'd163, 8'd166, 8'd172, 8'd184}, '{8'd179, 8'd167, 8'd173, 8'd185}, '{8'd171, 8'd182, 8'd174, 8'd186}, '{8'd187, 8'd183, 8'd175, 8'd187}, '{8'd167, 8'd174, 8'd188, 8'd188}, '{8'd183, 8'd175, 8'd189, 8'd189}, '{8'd175, 8'd190, 8'd190, 8'd190}, '{8'd191, 8'd191, 8'd191, 8'd191},
      '{8'd192, 8'd192, 8'd192, 8'd192}, '{8'd208, 8'd193, 8'd193, 8'd193}, '{8'd200, 8'd208, 8'd194, 8'd194}, '{8'd216, 8'd209, 8'd195, 8'd195}, '{8'd196, 8'd200, 8'd208, 8'd196}, '{8'd212, 8'd201, 8'd209, 8'd197}, '{8'd204, 8'd216, 8'd210, 8'd198}, '{8'd220, 8'd217, 8'd211, 8'd199},
      '{8'd193, 8'd194, 8'd196, 8'd200}, '{8'd209, 8'd195, 8'd197, 8'd201}, '{8'd201, 8'd210, 8'd198, 8'd202}, '{8'd217, 8'd211, 8'd199, 8'd203}, '{8'd197, 8'd202, 8'd212, 8'd204}, '{8'd213, 8'd203, 8'd213, 8'd205}, '{8'd205, 8'd218, 8'd214, 8'd206}, '{8'd221, 8'd219, 8'd215, 8'd207},
      '{8'd194, 8'd196, 8'd200, 8'd208}, '{8'd210, 8'd197, 8'd201, 8'd209}, '{8'd202, 8'd212, 8'd202, 8'd210}, '{8'd218, 8'd213, 8'd203, 8'd211}, '{8'd198, 8'd204, 8'd216, 8'd212}, '{8'd214, 8'd205, 8'd217, 8'd213}, '{8'd206, 8'd220, 8'd218, 8'd214}, '{8'd222, 8'd221, 8'd219, 8'd215},
      '{8'd195, 8'd198, 8'd204, 8'd216}, '{8'd211, 8'd199, 8'd205, 8'd217}, '{8'd203, 8'd214, 8'd206, 8'd218}, '{8'd219, 8'd215, 8'd207, 8'd219}, '{8'd199, 8'd206, 8'd220, 8'd220}, '{8'd215, 8'd207, 8'd221, 8'd221}, '{8'd207, 8'd222, 8'd222, 8'd222}, '{8'd223, 8'd223, 8'd223, 8'd223},
      '{8'd224, 8'd224, 8'd224, 8'd224}, '{8'd240, 8'd225, 8'd225, 8'd225}, '{8'd232, 8'd240, 8'd226, 8'd226}, '{8'd248, 8'd241, 8'd227, 8'd227}, '{8'd228, 8'd232, 8'd240, 8'd228}, '{8'd244, 8'd233, 8'd241, 8'd229}, '{8'd236, 8'd248, 8'd242, 8'd230}, '{8'd252, 8'd249, 8'd243, 8'd231},
      '{8'd225, 8'd226, 8'd228, 8'd232}, '{8'd241, 8'd227, 8'd229, 8'd233}, '{8'd233, 8'd242, 8'd230, 8'd234}, '{8'd249, 8'd243, 8'd231, 8'd235}, '{8'd229, 8'd234, 8'd244, 8'd236}, '{8'd245, 8'd235, 8'd245, 8'd237}, '{8'd237, 8'd250, 8'd246, 8'd238}, '{8'd253, 8'd251, 8'd247, 8'd239},
      '{8'd226, 8'd228, 8'd232, 8'd240}, '{8'd242, 8'd229, 8'd233, 8'd241}, '{8'd234, 8'd244, 8'd234, 8'd242}, '{8'd250, 8'd245, 8'd235, 8'd243}, '{8'd230, 8'd236, 8'd248, 8'd244}, '{8'd246, 8'd237, 8'd249, 8'd245}, '{8'd238, 8'd252, 8'd250, 8'd246}, '{8'd254, 8'd253, 8'd251, 8'd247},
      '{8'd227, 8'd230, 8'd236, 8'd248}, '{8'd243, 8'd231, 8'd237, 8'd249}, '{8'd235, 8'd246, 8'd238, 8'd250}, '{8'd251, 8'd247, 8'd239, 8'd251}, '{8'd231, 8'd238, 8'd252, 8'd252}, '{8'd247, 8'd239, 8'd253, 8'd253}, '{8'd239, 8'd254, 8'd254, 8'd254}, '{8'd255, 8'd255, 8'd255, 8'd255}
    };
    automatic logic [9-1:0] lut_16lane [0:511][0:3] = '{
      '{9'd000, 9'd000, 9'd000, 9'd000}, '{9'd016, 9'd001, 9'd001, 9'd001}, '{9'd008, 9'd016, 9'd002, 9'd002}, '{9'd024, 9'd017, 9'd003, 9'd003}, '{9'd004, 9'd008, 9'd016, 9'd004}, '{9'd020, 9'd009, 9'd017, 9'd005}, '{9'd012, 9'd024, 9'd018, 9'd006}, '{9'd028, 9'd025, 9'd019, 9'd007},
      '{9'd001, 9'd002, 9'd004, 9'd008}, '{9'd017, 9'd003, 9'd005, 9'd009}, '{9'd009, 9'd018, 9'd006, 9'd010}, '{9'd025, 9'd019, 9'd007, 9'd011}, '{9'd005, 9'd010, 9'd020, 9'd012}, '{9'd021, 9'd011, 9'd021, 9'd013}, '{9'd013, 9'd026, 9'd022, 9'd014}, '{9'd029, 9'd027, 9'd023, 9'd015},
      '{9'd002, 9'd004, 9'd008, 9'd016}, '{9'd018, 9'd005, 9'd009, 9'd017}, '{9'd010, 9'd020, 9'd010, 9'd018}, '{9'd026, 9'd021, 9'd011, 9'd019}, '{9'd006, 9'd012, 9'd024, 9'd020}, '{9'd022, 9'd013, 9'd025, 9'd021}, '{9'd014, 9'd028, 9'd026, 9'd022}, '{9'd030, 9'd029, 9'd027, 9'd023},
      '{9'd003, 9'd006, 9'd012, 9'd024}, '{9'd019, 9'd007, 9'd013, 9'd025}, '{9'd011, 9'd022, 9'd014, 9'd026}, '{9'd027, 9'd023, 9'd015, 9'd027}, '{9'd007, 9'd014, 9'd028, 9'd028}, '{9'd023, 9'd015, 9'd029, 9'd029}, '{9'd015, 9'd030, 9'd030, 9'd030}, '{9'd031, 9'd031, 9'd031, 9'd031},
      '{9'd032, 9'd032, 9'd032, 9'd032}, '{9'd048, 9'd033, 9'd033, 9'd033}, '{9'd040, 9'd048, 9'd034, 9'd034}, '{9'd056, 9'd049, 9'd035, 9'd035}, '{9'd036, 9'd040, 9'd048, 9'd036}, '{9'd052, 9'd041, 9'd049, 9'd037}, '{9'd044, 9'd056, 9'd050, 9'd038}, '{9'd060, 9'd057, 9'd051, 9'd039},
      '{9'd033, 9'd034, 9'd036, 9'd040}, '{9'd049, 9'd035, 9'd037, 9'd041}, '{9'd041, 9'd050, 9'd038, 9'd042}, '{9'd057, 9'd051, 9'd039, 9'd043}, '{9'd037, 9'd042, 9'd052, 9'd044}, '{9'd053, 9'd043, 9'd053, 9'd045}, '{9'd045, 9'd058, 9'd054, 9'd046}, '{9'd061, 9'd059, 9'd055, 9'd047},
      '{9'd034, 9'd036, 9'd040, 9'd048}, '{9'd050, 9'd037, 9'd041, 9'd049}, '{9'd042, 9'd052, 9'd042, 9'd050}, '{9'd058, 9'd053, 9'd043, 9'd051}, '{9'd038, 9'd044, 9'd056, 9'd052}, '{9'd054, 9'd045, 9'd057, 9'd053}, '{9'd046, 9'd060, 9'd058, 9'd054}, '{9'd062, 9'd061, 9'd059, 9'd055},
      '{9'd035, 9'd038, 9'd044, 9'd056}, '{9'd051, 9'd039, 9'd045, 9'd057}, '{9'd043, 9'd054, 9'd046, 9'd058}, '{9'd059, 9'd055, 9'd047, 9'd059}, '{9'd039, 9'd046, 9'd060, 9'd060}, '{9'd055, 9'd047, 9'd061, 9'd061}, '{9'd047, 9'd062, 9'd062, 9'd062}, '{9'd063, 9'd063, 9'd063, 9'd063},
      '{9'd064, 9'd064, 9'd064, 9'd064}, '{9'd080, 9'd065, 9'd065, 9'd065}, '{9'd072, 9'd080, 9'd066, 9'd066}, '{9'd088, 9'd081, 9'd067, 9'd067}, '{9'd068, 9'd072, 9'd080, 9'd068}, '{9'd084, 9'd073, 9'd081, 9'd069}, '{9'd076, 9'd088, 9'd082, 9'd070}, '{9'd092, 9'd089, 9'd083, 9'd071},
      '{9'd065, 9'd066, 9'd068, 9'd072}, '{9'd081, 9'd067, 9'd069, 9'd073}, '{9'd073, 9'd082, 9'd070, 9'd074}, '{9'd089, 9'd083, 9'd071, 9'd075}, '{9'd069, 9'd074, 9'd084, 9'd076}, '{9'd085, 9'd075, 9'd085, 9'd077}, '{9'd077, 9'd090, 9'd086, 9'd078}, '{9'd093, 9'd091, 9'd087, 9'd079},
      '{9'd066, 9'd068, 9'd072, 9'd080}, '{9'd082, 9'd069, 9'd073, 9'd081}, '{9'd074, 9'd084, 9'd074, 9'd082}, '{9'd090, 9'd085, 9'd075, 9'd083}, '{9'd070, 9'd076, 9'd088, 9'd084}, '{9'd086, 9'd077, 9'd089, 9'd085}, '{9'd078, 9'd092, 9'd090, 9'd086}, '{9'd094, 9'd093, 9'd091, 9'd087},
      '{9'd067, 9'd070, 9'd076, 9'd088}, '{9'd083, 9'd071, 9'd077, 9'd089}, '{9'd075, 9'd086, 9'd078, 9'd090}, '{9'd091, 9'd087, 9'd079, 9'd091}, '{9'd071, 9'd078, 9'd092, 9'd092}, '{9'd087, 9'd079, 9'd093, 9'd093}, '{9'd079, 9'd094, 9'd094, 9'd094}, '{9'd095, 9'd095, 9'd095, 9'd095},
      '{9'd096, 9'd096, 9'd096, 9'd096}, '{9'd112, 9'd097, 9'd097, 9'd097}, '{9'd104, 9'd112, 9'd098, 9'd098}, '{9'd120, 9'd113, 9'd099, 9'd099}, '{9'd100, 9'd104, 9'd112, 9'd100}, '{9'd116, 9'd105, 9'd113, 9'd101}, '{9'd108, 9'd120, 9'd114, 9'd102}, '{9'd124, 9'd121, 9'd115, 9'd103},
      '{9'd097, 9'd098, 9'd100, 9'd104}, '{9'd113, 9'd099, 9'd101, 9'd105}, '{9'd105, 9'd114, 9'd102, 9'd106}, '{9'd121, 9'd115, 9'd103, 9'd107}, '{9'd101, 9'd106, 9'd116, 9'd108}, '{9'd117, 9'd107, 9'd117, 9'd109}, '{9'd109, 9'd122, 9'd118, 9'd110}, '{9'd125, 9'd123, 9'd119, 9'd111},
      '{9'd098, 9'd100, 9'd104, 9'd112}, '{9'd114, 9'd101, 9'd105, 9'd113}, '{9'd106, 9'd116, 9'd106, 9'd114}, '{9'd122, 9'd117, 9'd107, 9'd115}, '{9'd102, 9'd108, 9'd120, 9'd116}, '{9'd118, 9'd109, 9'd121, 9'd117}, '{9'd110, 9'd124, 9'd122, 9'd118}, '{9'd126, 9'd125, 9'd123, 9'd119},
      '{9'd099, 9'd102, 9'd108, 9'd120}, '{9'd115, 9'd103, 9'd109, 9'd121}, '{9'd107, 9'd118, 9'd110, 9'd122}, '{9'd123, 9'd119, 9'd111, 9'd123}, '{9'd103, 9'd110, 9'd124, 9'd124}, '{9'd119, 9'd111, 9'd125, 9'd125}, '{9'd111, 9'd126, 9'd126, 9'd126}, '{9'd127, 9'd127, 9'd127, 9'd127},
      '{9'd128, 9'd128, 9'd128, 9'd128}, '{9'd144, 9'd129, 9'd129, 9'd129}, '{9'd136, 9'd144, 9'd130, 9'd130}, '{9'd152, 9'd145, 9'd131, 9'd131}, '{9'd132, 9'd136, 9'd144, 9'd132}, '{9'd148, 9'd137, 9'd145, 9'd133}, '{9'd140, 9'd152, 9'd146, 9'd134}, '{9'd156, 9'd153, 9'd147, 9'd135},
      '{9'd129, 9'd130, 9'd132, 9'd136}, '{9'd145, 9'd131, 9'd133, 9'd137}, '{9'd137, 9'd146, 9'd134, 9'd138}, '{9'd153, 9'd147, 9'd135, 9'd139}, '{9'd133, 9'd138, 9'd148, 9'd140}, '{9'd149, 9'd139, 9'd149, 9'd141}, '{9'd141, 9'd154, 9'd150, 9'd142}, '{9'd157, 9'd155, 9'd151, 9'd143},
      '{9'd130, 9'd132, 9'd136, 9'd144}, '{9'd146, 9'd133, 9'd137, 9'd145}, '{9'd138, 9'd148, 9'd138, 9'd146}, '{9'd154, 9'd149, 9'd139, 9'd147}, '{9'd134, 9'd140, 9'd152, 9'd148}, '{9'd150, 9'd141, 9'd153, 9'd149}, '{9'd142, 9'd156, 9'd154, 9'd150}, '{9'd158, 9'd157, 9'd155, 9'd151},
      '{9'd131, 9'd134, 9'd140, 9'd152}, '{9'd147, 9'd135, 9'd141, 9'd153}, '{9'd139, 9'd150, 9'd142, 9'd154}, '{9'd155, 9'd151, 9'd143, 9'd155}, '{9'd135, 9'd142, 9'd156, 9'd156}, '{9'd151, 9'd143, 9'd157, 9'd157}, '{9'd143, 9'd158, 9'd158, 9'd158}, '{9'd159, 9'd159, 9'd159, 9'd159},
      '{9'd160, 9'd160, 9'd160, 9'd160}, '{9'd176, 9'd161, 9'd161, 9'd161}, '{9'd168, 9'd176, 9'd162, 9'd162}, '{9'd184, 9'd177, 9'd163, 9'd163}, '{9'd164, 9'd168, 9'd176, 9'd164}, '{9'd180, 9'd169, 9'd177, 9'd165}, '{9'd172, 9'd184, 9'd178, 9'd166}, '{9'd188, 9'd185, 9'd179, 9'd167},
      '{9'd161, 9'd162, 9'd164, 9'd168}, '{9'd177, 9'd163, 9'd165, 9'd169}, '{9'd169, 9'd178, 9'd166, 9'd170}, '{9'd185, 9'd179, 9'd167, 9'd171}, '{9'd165, 9'd170, 9'd180, 9'd172}, '{9'd181, 9'd171, 9'd181, 9'd173}, '{9'd173, 9'd186, 9'd182, 9'd174}, '{9'd189, 9'd187, 9'd183, 9'd175},
      '{9'd162, 9'd164, 9'd168, 9'd176}, '{9'd178, 9'd165, 9'd169, 9'd177}, '{9'd170, 9'd180, 9'd170, 9'd178}, '{9'd186, 9'd181, 9'd171, 9'd179}, '{9'd166, 9'd172, 9'd184, 9'd180}, '{9'd182, 9'd173, 9'd185, 9'd181}, '{9'd174, 9'd188, 9'd186, 9'd182}, '{9'd190, 9'd189, 9'd187, 9'd183},
      '{9'd163, 9'd166, 9'd172, 9'd184}, '{9'd179, 9'd167, 9'd173, 9'd185}, '{9'd171, 9'd182, 9'd174, 9'd186}, '{9'd187, 9'd183, 9'd175, 9'd187}, '{9'd167, 9'd174, 9'd188, 9'd188}, '{9'd183, 9'd175, 9'd189, 9'd189}, '{9'd175, 9'd190, 9'd190, 9'd190}, '{9'd191, 9'd191, 9'd191, 9'd191},
      '{9'd192, 9'd192, 9'd192, 9'd192}, '{9'd208, 9'd193, 9'd193, 9'd193}, '{9'd200, 9'd208, 9'd194, 9'd194}, '{9'd216, 9'd209, 9'd195, 9'd195}, '{9'd196, 9'd200, 9'd208, 9'd196}, '{9'd212, 9'd201, 9'd209, 9'd197}, '{9'd204, 9'd216, 9'd210, 9'd198}, '{9'd220, 9'd217, 9'd211, 9'd199},
      '{9'd193, 9'd194, 9'd196, 9'd200}, '{9'd209, 9'd195, 9'd197, 9'd201}, '{9'd201, 9'd210, 9'd198, 9'd202}, '{9'd217, 9'd211, 9'd199, 9'd203}, '{9'd197, 9'd202, 9'd212, 9'd204}, '{9'd213, 9'd203, 9'd213, 9'd205}, '{9'd205, 9'd218, 9'd214, 9'd206}, '{9'd221, 9'd219, 9'd215, 9'd207},
      '{9'd194, 9'd196, 9'd200, 9'd208}, '{9'd210, 9'd197, 9'd201, 9'd209}, '{9'd202, 9'd212, 9'd202, 9'd210}, '{9'd218, 9'd213, 9'd203, 9'd211}, '{9'd198, 9'd204, 9'd216, 9'd212}, '{9'd214, 9'd205, 9'd217, 9'd213}, '{9'd206, 9'd220, 9'd218, 9'd214}, '{9'd222, 9'd221, 9'd219, 9'd215},
      '{9'd195, 9'd198, 9'd204, 9'd216}, '{9'd211, 9'd199, 9'd205, 9'd217}, '{9'd203, 9'd214, 9'd206, 9'd218}, '{9'd219, 9'd215, 9'd207, 9'd219}, '{9'd199, 9'd206, 9'd220, 9'd220}, '{9'd215, 9'd207, 9'd221, 9'd221}, '{9'd207, 9'd222, 9'd222, 9'd222}, '{9'd223, 9'd223, 9'd223, 9'd223},
      '{9'd224, 9'd224, 9'd224, 9'd224}, '{9'd240, 9'd225, 9'd225, 9'd225}, '{9'd232, 9'd240, 9'd226, 9'd226}, '{9'd248, 9'd241, 9'd227, 9'd227}, '{9'd228, 9'd232, 9'd240, 9'd228}, '{9'd244, 9'd233, 9'd241, 9'd229}, '{9'd236, 9'd248, 9'd242, 9'd230}, '{9'd252, 9'd249, 9'd243, 9'd231},
      '{9'd225, 9'd226, 9'd228, 9'd232}, '{9'd241, 9'd227, 9'd229, 9'd233}, '{9'd233, 9'd242, 9'd230, 9'd234}, '{9'd249, 9'd243, 9'd231, 9'd235}, '{9'd229, 9'd234, 9'd244, 9'd236}, '{9'd245, 9'd235, 9'd245, 9'd237}, '{9'd237, 9'd250, 9'd246, 9'd238}, '{9'd253, 9'd251, 9'd247, 9'd239},
      '{9'd226, 9'd228, 9'd232, 9'd240}, '{9'd242, 9'd229, 9'd233, 9'd241}, '{9'd234, 9'd244, 9'd234, 9'd242}, '{9'd250, 9'd245, 9'd235, 9'd243}, '{9'd230, 9'd236, 9'd248, 9'd244}, '{9'd246, 9'd237, 9'd249, 9'd245}, '{9'd238, 9'd252, 9'd250, 9'd246}, '{9'd254, 9'd253, 9'd251, 9'd247},
      '{9'd227, 9'd230, 9'd236, 9'd248}, '{9'd243, 9'd231, 9'd237, 9'd249}, '{9'd235, 9'd246, 9'd238, 9'd250}, '{9'd251, 9'd247, 9'd239, 9'd251}, '{9'd231, 9'd238, 9'd252, 9'd252}, '{9'd247, 9'd239, 9'd253, 9'd253}, '{9'd239, 9'd254, 9'd254, 9'd254}, '{9'd255, 9'd255, 9'd255, 9'd255},
      '{9'd256, 9'd256, 9'd256, 9'd256}, '{9'd272, 9'd257, 9'd257, 9'd257}, '{9'd264, 9'd272, 9'd258, 9'd258}, '{9'd280, 9'd273, 9'd259, 9'd259}, '{9'd260, 9'd264, 9'd272, 9'd260}, '{9'd276, 9'd265, 9'd273, 9'd261}, '{9'd268, 9'd280, 9'd274, 9'd262}, '{9'd284, 9'd281, 9'd275, 9'd263},
      '{9'd257, 9'd258, 9'd260, 9'd264}, '{9'd273, 9'd259, 9'd261, 9'd265}, '{9'd265, 9'd274, 9'd262, 9'd266}, '{9'd281, 9'd275, 9'd263, 9'd267}, '{9'd261, 9'd266, 9'd276, 9'd268}, '{9'd277, 9'd267, 9'd277, 9'd269}, '{9'd269, 9'd282, 9'd278, 9'd270}, '{9'd285, 9'd283, 9'd279, 9'd271},
      '{9'd258, 9'd260, 9'd264, 9'd272}, '{9'd274, 9'd261, 9'd265, 9'd273}, '{9'd266, 9'd276, 9'd266, 9'd274}, '{9'd282, 9'd277, 9'd267, 9'd275}, '{9'd262, 9'd268, 9'd280, 9'd276}, '{9'd278, 9'd269, 9'd281, 9'd277}, '{9'd270, 9'd284, 9'd282, 9'd278}, '{9'd286, 9'd285, 9'd283, 9'd279},
      '{9'd259, 9'd262, 9'd268, 9'd280}, '{9'd275, 9'd263, 9'd269, 9'd281}, '{9'd267, 9'd278, 9'd270, 9'd282}, '{9'd283, 9'd279, 9'd271, 9'd283}, '{9'd263, 9'd270, 9'd284, 9'd284}, '{9'd279, 9'd271, 9'd285, 9'd285}, '{9'd271, 9'd286, 9'd286, 9'd286}, '{9'd287, 9'd287, 9'd287, 9'd287},
      '{9'd288, 9'd288, 9'd288, 9'd288}, '{9'd304, 9'd289, 9'd289, 9'd289}, '{9'd296, 9'd304, 9'd290, 9'd290}, '{9'd312, 9'd305, 9'd291, 9'd291}, '{9'd292, 9'd296, 9'd304, 9'd292}, '{9'd308, 9'd297, 9'd305, 9'd293}, '{9'd300, 9'd312, 9'd306, 9'd294}, '{9'd316, 9'd313, 9'd307, 9'd295},
      '{9'd289, 9'd290, 9'd292, 9'd296}, '{9'd305, 9'd291, 9'd293, 9'd297}, '{9'd297, 9'd306, 9'd294, 9'd298}, '{9'd313, 9'd307, 9'd295, 9'd299}, '{9'd293, 9'd298, 9'd308, 9'd300}, '{9'd309, 9'd299, 9'd309, 9'd301}, '{9'd301, 9'd314, 9'd310, 9'd302}, '{9'd317, 9'd315, 9'd311, 9'd303},
      '{9'd290, 9'd292, 9'd296, 9'd304}, '{9'd306, 9'd293, 9'd297, 9'd305}, '{9'd298, 9'd308, 9'd298, 9'd306}, '{9'd314, 9'd309, 9'd299, 9'd307}, '{9'd294, 9'd300, 9'd312, 9'd308}, '{9'd310, 9'd301, 9'd313, 9'd309}, '{9'd302, 9'd316, 9'd314, 9'd310}, '{9'd318, 9'd317, 9'd315, 9'd311},
      '{9'd291, 9'd294, 9'd300, 9'd312}, '{9'd307, 9'd295, 9'd301, 9'd313}, '{9'd299, 9'd310, 9'd302, 9'd314}, '{9'd315, 9'd311, 9'd303, 9'd315}, '{9'd295, 9'd302, 9'd316, 9'd316}, '{9'd311, 9'd303, 9'd317, 9'd317}, '{9'd303, 9'd318, 9'd318, 9'd318}, '{9'd319, 9'd319, 9'd319, 9'd319},
      '{9'd320, 9'd320, 9'd320, 9'd320}, '{9'd336, 9'd321, 9'd321, 9'd321}, '{9'd328, 9'd336, 9'd322, 9'd322}, '{9'd344, 9'd337, 9'd323, 9'd323}, '{9'd324, 9'd328, 9'd336, 9'd324}, '{9'd340, 9'd329, 9'd337, 9'd325}, '{9'd332, 9'd344, 9'd338, 9'd326}, '{9'd348, 9'd345, 9'd339, 9'd327},
      '{9'd321, 9'd322, 9'd324, 9'd328}, '{9'd337, 9'd323, 9'd325, 9'd329}, '{9'd329, 9'd338, 9'd326, 9'd330}, '{9'd345, 9'd339, 9'd327, 9'd331}, '{9'd325, 9'd330, 9'd340, 9'd332}, '{9'd341, 9'd331, 9'd341, 9'd333}, '{9'd333, 9'd346, 9'd342, 9'd334}, '{9'd349, 9'd347, 9'd343, 9'd335},
      '{9'd322, 9'd324, 9'd328, 9'd336}, '{9'd338, 9'd325, 9'd329, 9'd337}, '{9'd330, 9'd340, 9'd330, 9'd338}, '{9'd346, 9'd341, 9'd331, 9'd339}, '{9'd326, 9'd332, 9'd344, 9'd340}, '{9'd342, 9'd333, 9'd345, 9'd341}, '{9'd334, 9'd348, 9'd346, 9'd342}, '{9'd350, 9'd349, 9'd347, 9'd343},
      '{9'd323, 9'd326, 9'd332, 9'd344}, '{9'd339, 9'd327, 9'd333, 9'd345}, '{9'd331, 9'd342, 9'd334, 9'd346}, '{9'd347, 9'd343, 9'd335, 9'd347}, '{9'd327, 9'd334, 9'd348, 9'd348}, '{9'd343, 9'd335, 9'd349, 9'd349}, '{9'd335, 9'd350, 9'd350, 9'd350}, '{9'd351, 9'd351, 9'd351, 9'd351},
      '{9'd352, 9'd352, 9'd352, 9'd352}, '{9'd368, 9'd353, 9'd353, 9'd353}, '{9'd360, 9'd368, 9'd354, 9'd354}, '{9'd376, 9'd369, 9'd355, 9'd355}, '{9'd356, 9'd360, 9'd368, 9'd356}, '{9'd372, 9'd361, 9'd369, 9'd357}, '{9'd364, 9'd376, 9'd370, 9'd358}, '{9'd380, 9'd377, 9'd371, 9'd359},
      '{9'd353, 9'd354, 9'd356, 9'd360}, '{9'd369, 9'd355, 9'd357, 9'd361}, '{9'd361, 9'd370, 9'd358, 9'd362}, '{9'd377, 9'd371, 9'd359, 9'd363}, '{9'd357, 9'd362, 9'd372, 9'd364}, '{9'd373, 9'd363, 9'd373, 9'd365}, '{9'd365, 9'd378, 9'd374, 9'd366}, '{9'd381, 9'd379, 9'd375, 9'd367},
      '{9'd354, 9'd356, 9'd360, 9'd368}, '{9'd370, 9'd357, 9'd361, 9'd369}, '{9'd362, 9'd372, 9'd362, 9'd370}, '{9'd378, 9'd373, 9'd363, 9'd371}, '{9'd358, 9'd364, 9'd376, 9'd372}, '{9'd374, 9'd365, 9'd377, 9'd373}, '{9'd366, 9'd380, 9'd378, 9'd374}, '{9'd382, 9'd381, 9'd379, 9'd375},
      '{9'd355, 9'd358, 9'd364, 9'd376}, '{9'd371, 9'd359, 9'd365, 9'd377}, '{9'd363, 9'd374, 9'd366, 9'd378}, '{9'd379, 9'd375, 9'd367, 9'd379}, '{9'd359, 9'd366, 9'd380, 9'd380}, '{9'd375, 9'd367, 9'd381, 9'd381}, '{9'd367, 9'd382, 9'd382, 9'd382}, '{9'd383, 9'd383, 9'd383, 9'd383},
      '{9'd384, 9'd384, 9'd384, 9'd384}, '{9'd400, 9'd385, 9'd385, 9'd385}, '{9'd392, 9'd400, 9'd386, 9'd386}, '{9'd408, 9'd401, 9'd387, 9'd387}, '{9'd388, 9'd392, 9'd400, 9'd388}, '{9'd404, 9'd393, 9'd401, 9'd389}, '{9'd396, 9'd408, 9'd402, 9'd390}, '{9'd412, 9'd409, 9'd403, 9'd391},
      '{9'd385, 9'd386, 9'd388, 9'd392}, '{9'd401, 9'd387, 9'd389, 9'd393}, '{9'd393, 9'd402, 9'd390, 9'd394}, '{9'd409, 9'd403, 9'd391, 9'd395}, '{9'd389, 9'd394, 9'd404, 9'd396}, '{9'd405, 9'd395, 9'd405, 9'd397}, '{9'd397, 9'd410, 9'd406, 9'd398}, '{9'd413, 9'd411, 9'd407, 9'd399},
      '{9'd386, 9'd388, 9'd392, 9'd400}, '{9'd402, 9'd389, 9'd393, 9'd401}, '{9'd394, 9'd404, 9'd394, 9'd402}, '{9'd410, 9'd405, 9'd395, 9'd403}, '{9'd390, 9'd396, 9'd408, 9'd404}, '{9'd406, 9'd397, 9'd409, 9'd405}, '{9'd398, 9'd412, 9'd410, 9'd406}, '{9'd414, 9'd413, 9'd411, 9'd407},
      '{9'd387, 9'd390, 9'd396, 9'd408}, '{9'd403, 9'd391, 9'd397, 9'd409}, '{9'd395, 9'd406, 9'd398, 9'd410}, '{9'd411, 9'd407, 9'd399, 9'd411}, '{9'd391, 9'd398, 9'd412, 9'd412}, '{9'd407, 9'd399, 9'd413, 9'd413}, '{9'd399, 9'd414, 9'd414, 9'd414}, '{9'd415, 9'd415, 9'd415, 9'd415},
      '{9'd416, 9'd416, 9'd416, 9'd416}, '{9'd432, 9'd417, 9'd417, 9'd417}, '{9'd424, 9'd432, 9'd418, 9'd418}, '{9'd440, 9'd433, 9'd419, 9'd419}, '{9'd420, 9'd424, 9'd432, 9'd420}, '{9'd436, 9'd425, 9'd433, 9'd421}, '{9'd428, 9'd440, 9'd434, 9'd422}, '{9'd444, 9'd441, 9'd435, 9'd423},
      '{9'd417, 9'd418, 9'd420, 9'd424}, '{9'd433, 9'd419, 9'd421, 9'd425}, '{9'd425, 9'd434, 9'd422, 9'd426}, '{9'd441, 9'd435, 9'd423, 9'd427}, '{9'd421, 9'd426, 9'd436, 9'd428}, '{9'd437, 9'd427, 9'd437, 9'd429}, '{9'd429, 9'd442, 9'd438, 9'd430}, '{9'd445, 9'd443, 9'd439, 9'd431},
      '{9'd418, 9'd420, 9'd424, 9'd432}, '{9'd434, 9'd421, 9'd425, 9'd433}, '{9'd426, 9'd436, 9'd426, 9'd434}, '{9'd442, 9'd437, 9'd427, 9'd435}, '{9'd422, 9'd428, 9'd440, 9'd436}, '{9'd438, 9'd429, 9'd441, 9'd437}, '{9'd430, 9'd444, 9'd442, 9'd438}, '{9'd446, 9'd445, 9'd443, 9'd439},
      '{9'd419, 9'd422, 9'd428, 9'd440}, '{9'd435, 9'd423, 9'd429, 9'd441}, '{9'd427, 9'd438, 9'd430, 9'd442}, '{9'd443, 9'd439, 9'd431, 9'd443}, '{9'd423, 9'd430, 9'd444, 9'd444}, '{9'd439, 9'd431, 9'd445, 9'd445}, '{9'd431, 9'd446, 9'd446, 9'd446}, '{9'd447, 9'd447, 9'd447, 9'd447},
      '{9'd448, 9'd448, 9'd448, 9'd448}, '{9'd464, 9'd449, 9'd449, 9'd449}, '{9'd456, 9'd464, 9'd450, 9'd450}, '{9'd472, 9'd465, 9'd451, 9'd451}, '{9'd452, 9'd456, 9'd464, 9'd452}, '{9'd468, 9'd457, 9'd465, 9'd453}, '{9'd460, 9'd472, 9'd466, 9'd454}, '{9'd476, 9'd473, 9'd467, 9'd455},
      '{9'd449, 9'd450, 9'd452, 9'd456}, '{9'd465, 9'd451, 9'd453, 9'd457}, '{9'd457, 9'd466, 9'd454, 9'd458}, '{9'd473, 9'd467, 9'd455, 9'd459}, '{9'd453, 9'd458, 9'd468, 9'd460}, '{9'd469, 9'd459, 9'd469, 9'd461}, '{9'd461, 9'd474, 9'd470, 9'd462}, '{9'd477, 9'd475, 9'd471, 9'd463},
      '{9'd450, 9'd452, 9'd456, 9'd464}, '{9'd466, 9'd453, 9'd457, 9'd465}, '{9'd458, 9'd468, 9'd458, 9'd466}, '{9'd474, 9'd469, 9'd459, 9'd467}, '{9'd454, 9'd460, 9'd472, 9'd468}, '{9'd470, 9'd461, 9'd473, 9'd469}, '{9'd462, 9'd476, 9'd474, 9'd470}, '{9'd478, 9'd477, 9'd475, 9'd471},
      '{9'd451, 9'd454, 9'd460, 9'd472}, '{9'd467, 9'd455, 9'd461, 9'd473}, '{9'd459, 9'd470, 9'd462, 9'd474}, '{9'd475, 9'd471, 9'd463, 9'd475}, '{9'd455, 9'd462, 9'd476, 9'd476}, '{9'd471, 9'd463, 9'd477, 9'd477}, '{9'd463, 9'd478, 9'd478, 9'd478}, '{9'd479, 9'd479, 9'd479, 9'd479},
      '{9'd480, 9'd480, 9'd480, 9'd480}, '{9'd496, 9'd481, 9'd481, 9'd481}, '{9'd488, 9'd496, 9'd482, 9'd482}, '{9'd504, 9'd497, 9'd483, 9'd483}, '{9'd484, 9'd488, 9'd496, 9'd484}, '{9'd500, 9'd489, 9'd497, 9'd485}, '{9'd492, 9'd504, 9'd498, 9'd486}, '{9'd508, 9'd505, 9'd499, 9'd487},
      '{9'd481, 9'd482, 9'd484, 9'd488}, '{9'd497, 9'd483, 9'd485, 9'd489}, '{9'd489, 9'd498, 9'd486, 9'd490}, '{9'd505, 9'd499, 9'd487, 9'd491}, '{9'd485, 9'd490, 9'd500, 9'd492}, '{9'd501, 9'd491, 9'd501, 9'd493}, '{9'd493, 9'd506, 9'd502, 9'd494}, '{9'd509, 9'd507, 9'd503, 9'd495},
      '{9'd482, 9'd484, 9'd488, 9'd496}, '{9'd498, 9'd485, 9'd489, 9'd497}, '{9'd490, 9'd500, 9'd490, 9'd498}, '{9'd506, 9'd501, 9'd491, 9'd499}, '{9'd486, 9'd492, 9'd504, 9'd500}, '{9'd502, 9'd493, 9'd505, 9'd501}, '{9'd494, 9'd508, 9'd506, 9'd502}, '{9'd510, 9'd509, 9'd507, 9'd503},
      '{9'd483, 9'd486, 9'd492, 9'd504}, '{9'd499, 9'd487, 9'd493, 9'd505}, '{9'd491, 9'd502, 9'd494, 9'd506}, '{9'd507, 9'd503, 9'd495, 9'd507}, '{9'd487, 9'd494, 9'd508, 9'd508}, '{9'd503, 9'd495, 9'd509, 9'd509}, '{9'd495, 9'd510, 9'd510, 9'd510}, '{9'd511, 9'd511, 9'd511, 9'd511}
    };

    unique case (NrLanes)
      1 : return lut_1lane [shfNbIdx][ew];
      2 : return lut_2lane [shfNbIdx][ew];
      4 : return lut_4lane [shfNbIdx][ew];
      8 : return lut_8lane [shfNbIdx][ew];
      16: return lut_16lane[shfNbIdx][ew];
      default: return 0;
	  endcase
  endfunction

  // // Input shuffle index, output sequential index  
  // // Used in Shuffle Unit to convert shuffle index to sequential index
  // function automatic logic [{$clog2(riva_pkg::DLEN*riva_pkg::MaxNrLanes/4)}-1:0] query_seq_idx(input int NrLanes, input int shfNbIdx, input riscv_mv_pkg::vew_e ew);
  //   unique case (NrLanes)
  //     1: begin
  //       automatic logic [5-1:0] idx [0:3];
  //       for (int seqIdx = 0; seqIdx < 32; seqIdx++)
  //           idx[query_shf_idx(NrLanes, seqIdx, ew)] = seqIdx;
  //       return idx[shfNbIdx];
  //     end
  //     2: begin
  //       automatic logic [6-1:0] idx [0:3];
  //       for (int seqIdx = 0; seqIdx < 64; seqIdx++)
  //         idx[query_shf_idx(NrLanes, seqIdx, ew)] = seqIdx;
  //       return idx[shfNbIdx];
  //     end
  //     4: begin
  //       automatic logic [7-1:0] idx [0:3];
  //       for (int unsigned seqIdx = 0; seqIdx < 128; seqIdx++) begin
  //         automatic int unsigned shf_idx = query_shf_idx(NrLanes, seqIdx, ew);
  //         idx[shf_idx] = seqIdx;
  //         $display("idx[%0d] = %0d", shf_idx, seqIdx);
  //       end
  //       // print full idx
  //       for (int i = 0; i < 128; i++) begin
  //         $display("idx[%0d] = %0d", i, idx[i]);
  //       end
  //       return idx[shfNbIdx];
  //     end
  //     8: begin
  //       automatic logic [8-1:0] idx [0:3];
  //       for (int seqIdx = 0; seqIdx < 256; seqIdx++)
  //         idx[query_shf_idx(NrLanes, seqIdx, ew)] = seqIdx;
  //       return idx[shfNbIdx];
  //     end
  //     16: begin
  //       automatic logic [9-1:0] idx [0:3];
  //       for (int seqIdx = 0; seqIdx < 512; seqIdx++)
  //         idx[query_shf_idx(NrLanes, seqIdx, ew)] = seqIdx;
  //       return idx[shfNbIdx];
  //     end
  //     default: return 0;
  //   endcase
  // endfunction: query_seq_idx

  // // Input shuffle index, output sequential index for 2D column-major mode
  // // Used in Shuffle Unit to convert shuffle index to sequential index
  // function automatic logic [{$clog2(riva_pkg::DLEN*riva_pkg::MaxNrLanes/4)}-1:0] query_seq_idx_2d_cln(input int NrLanes, input int shfNbIdx, input riscv_mv_pkg::vew_e ew);
  //   unique case (NrLanes)
  //     1: begin
  //       automatic logic [5-1:0] idx [0:3];
  //       for (int seqIdx = 0; seqIdx < 32; seqIdx++)
  //           idx[query_shf_idx_2d_cln(NrLanes, seqIdx, ew)] = seqIdx;
  //       return idx[shfNbIdx];
  //     end
  //     2: begin
  //       automatic logic [6-1:0] idx [0:3];
  //       for (int seqIdx = 0; seqIdx < 64; seqIdx++)
  //         idx[query_shf_idx_2d_cln(NrLanes, seqIdx, ew)] = seqIdx;
  //       return idx[shfNbIdx];
  //     end
  //     4: begin
  //       automatic logic [7-1:0] idx [0:3];
  //       for (int seqIdx = 0; seqIdx < 128; seqIdx++)
  //         idx[query_shf_idx_2d_cln(NrLanes, seqIdx, ew)] = seqIdx;
  //       for (int i = 0; i < 4; i++) begin
  //          $display("idx[%0d] = %0d", i, idx[i]);
  //       end
  //       return idx[shfNbIdx];
  //     end
  //     8: begin
  //       automatic logic [8-1:0] idx [0:3];
  //       for (int seqIdx = 0; seqIdx < 256; seqIdx++)
  //         idx[query_shf_idx_2d_cln(NrLanes, seqIdx, ew)] = seqIdx;
  //       return idx[shfNbIdx];
  //     end
  //     16: begin
  //       automatic logic [9-1:0] idx [0:3];
  //       for (int seqIdx = 0; seqIdx < 512; seqIdx++)
  //         idx[query_shf_idx_2d_cln(NrLanes, seqIdx, ew)] = seqIdx;
  //       return idx[shfNbIdx];
  //     end
  //     default: return 0;
	//   endcase
  // endfunction: query_seq_idx_2d_cln

endpackage